------------------------------------------------------------
--author: tretterch
--date:	  03-15-2017
--Descr.: Implementation of cordic implementation for 
--	  exponential function
------------------------------------------------------------
--Rev	 author		date		comment
--0.1	tretterch     03-15-2017      initial implementation
------------------------------------------------------------

architecture RTL of Cordic is

begin

end architecture RTL
