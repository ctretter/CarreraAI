-- megafunction wizard: %ALTFP_EXP%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_EXP 

-- ============================================================
-- File Name: ALTFP_EXa.vhd
-- Megafunction Name(s):
-- 			ALTFP_EXP
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.0.0 Build 211 04/27/2016 SJ Standard Edition
-- ************************************************************


--Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altfp_exp CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=25 ROUNDING="TO_NEAREST" WIDTH_EXP=11 WIDTH_MAN=52 aclr clock data result
--VERSION_BEGIN 16.0 cbx_altfp_exp 2016:04:27:18:05:34:SJ cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_clshift 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_lpm_mux 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END


--altmult_opt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" LPM_PIPELINE=4 LPM_WIDTHA=60 LPM_WIDTHB=60 LPM_WIDTHP=120 aclr clken clock dataa datab result
--VERSION_BEGIN 16.0 cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END


--altmult_opt_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=90 aclr clken clock dataa datab result
--VERSION_BEGIN 16.0 cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altmult_opt_csa_ksf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (89 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (89 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (89 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altmult_opt_csa_ksf;

 ARCHITECTURE RTL OF ALTFP_EXa_altmult_opt_csa_ksf IS

	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub1_result;
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 90
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub1_result
	  );

 END RTL; --ALTFP_EXa_altmult_opt_csa_ksf

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 lpm_mult 3 reg 422 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altmult_opt_v4e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (59 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (59 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (119 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altmult_opt_v4e;

 ARCHITECTURE RTL OF ALTFP_EXa_altmult_opt_v4e IS

	 SIGNAL  wire_sum_result	:	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL	 car_two_adj_reg0	:	STD_LOGIC_VECTOR(89 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg0	:	STD_LOGIC_VECTOR(29 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg1	:	STD_LOGIC_VECTOR(29 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lsb_prod_wi_reg0	:	STD_LOGIC_VECTOR(59 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mid_prod_wi_reg0	:	STD_LOGIC_VECTOR(61 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 msb_prod_wi_reg0	:	STD_LOGIC_VECTOR(59 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sum_two_reg0	:	STD_LOGIC_VECTOR(89 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_compress_a_cout	:	STD_LOGIC;
	 SIGNAL  wire_compress_a_result	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_compress_b_cout	:	STD_LOGIC;
	 SIGNAL  wire_compress_b_result	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_lsb_prod_result	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_mid_prod_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_mid_prod_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_mid_prod_result	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_msb_prod_result	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4183w4192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4123w4293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4117w4303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4111w4313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4105w4323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4099w4333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4093w4343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4087w4353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4081w4363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4075w4373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4069w4383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4177w4203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4063w4393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4057w4403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4051w4413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4045w4423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4039w4433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4033w4443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4027w4453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4021w4463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4015w4473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4009w4483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4171w4213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4003w4493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3997w4503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3991w4513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3985w4523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3979w4533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3973w4543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3967w4553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3961w4563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3955w4573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3949w4583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4165w4223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3943w4593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3937w4603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3931w4613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3925w4623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3919w4633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3913w4643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3907w4653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3901w4663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3895w4673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3889w4683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4159w4233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3883w4693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3877w4703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3871w4713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3865w4723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3859w4733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3853w4743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3847w4753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3841w4763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3835w4773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3829w4783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4153w4243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3823w4793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3819w4803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3815w4813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3811w4823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3807w4833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3803w4843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3799w4853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3795w4863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3791w4873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3787w4883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4147w4253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3783w4893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3779w4903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3775w4913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3771w4923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3767w4933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3763w4943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3759w4953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3755w4963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3751w4973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3747w4983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4141w4263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3743w4993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3739w5003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3735w5013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3731w5023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3727w5033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3723w5043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3719w5053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3715w5063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3711w5073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range3705w5083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4135w4273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_neg_msb_range4129w4283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4190w5099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4292w5210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4302w5221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4312w5232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4322w5243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4332w5254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4342w5265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4352w5276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4362w5287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4372w5298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4382w5309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4202w5111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4392w5320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4402w5331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4412w5342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4422w5353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4432w5364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4442w5375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4452w5386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4462w5397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4472w5408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4482w5419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4212w5122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4492w5430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4502w5441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4512w5452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4522w5463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4532w5474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4542w5485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4552w5496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4562w5507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4572w5518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4582w5529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4222w5133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4592w5540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4602w5551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4612w5562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4622w5573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4632w5584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4642w5595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4652w5606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4662w5617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4672w5628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4682w5639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4232w5144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4692w5650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4702w5661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4712w5672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4722w5683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4732w5694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4742w5705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4752w5716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4762w5727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4772w5738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4782w5749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4242w5155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4792w5760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4802w5771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4812w5782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4822w5793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4832w5804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4842w5815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4852w5826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4862w5837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4872w5848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4882w5859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4252w5166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4892w5870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4902w5881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4912w5892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4922w5903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4932w5914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4942w5925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4952w5936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4962w5947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4972w5958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4982w5969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4262w5177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4992w5980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5002w5991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5012w6002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5022w6013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5032w6024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5042w6035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5052w6046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5062w6057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5072w6068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range5082w6079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4272w5188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_sum_one_range4282w5199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5094w5100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5094w5101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5206w5211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5206w5212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5217w5222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5217w5223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5228w5233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5228w5234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5239w5244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5239w5245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5250w5255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5250w5256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5261w5266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5261w5267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5272w5277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5272w5278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5283w5288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5283w5289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5294w5299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5294w5300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5305w5310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5305w5311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5107w5112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5107w5113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5316w5321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5316w5322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5327w5332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5327w5333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5338w5343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5338w5344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5349w5354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5349w5355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5360w5365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5360w5366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5371w5376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5371w5377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5382w5387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5382w5388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5393w5398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5393w5399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5404w5409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5404w5410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5415w5420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5415w5421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5118w5123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5118w5124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5426w5431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5426w5432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5437w5442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5437w5443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5448w5453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5448w5454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5459w5464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5459w5465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5470w5475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5470w5476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5481w5486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5481w5487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5492w5497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5492w5498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5503w5508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5503w5509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5514w5519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5514w5520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5525w5530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5525w5531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5129w5134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5129w5135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5536w5541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5536w5542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5547w5552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5547w5553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5558w5563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5558w5564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5569w5574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5569w5575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5580w5585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5580w5586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5591w5596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5591w5597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5602w5607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5602w5608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5613w5618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5613w5619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5624w5629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5624w5630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5635w5640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5635w5641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5140w5145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5140w5146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5646w5651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5646w5652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5657w5662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5657w5663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5668w5673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5668w5674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5679w5684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5679w5685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5690w5695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5690w5696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5701w5706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5701w5707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5712w5717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5712w5718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5723w5728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5723w5729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5734w5739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5734w5740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5745w5750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5745w5751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5151w5156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5151w5157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5756w5761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5756w5762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5767w5772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5767w5773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5778w5783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5778w5784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5789w5794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5789w5795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5800w5805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5800w5806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5811w5816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5811w5817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5822w5827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5822w5828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5833w5838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5833w5839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5844w5849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5844w5850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5855w5860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5855w5861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5162w5167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5162w5168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5866w5871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5866w5872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5877w5882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5877w5883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5888w5893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5888w5894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5899w5904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5899w5905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5910w5915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5910w5916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5921w5926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5921w5927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5932w5937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5932w5938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5943w5948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5943w5949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5954w5959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5954w5960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5965w5970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5965w5971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5173w5178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5173w5179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5976w5981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5976w5982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5987w5992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5987w5993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5998w6003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5998w6004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6009w6014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6009w6015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6020w6025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6020w6026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6031w6036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6031w6037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6042w6047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6042w6048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6053w6058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6053w6059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6064w6069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6064w6070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6075w6080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6075w6081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5184w5189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5184w5190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5195w5200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5195w5201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4187w4193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4187w4194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4289w4294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4289w4295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4299w4304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4299w4305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4309w4314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4309w4315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4319w4324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4319w4325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4329w4334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4329w4335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4339w4344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4339w4345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4349w4354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4349w4355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4359w4364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4359w4365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4369w4374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4369w4375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4379w4384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4379w4385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4199w4204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4199w4205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4389w4394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4389w4395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4399w4404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4399w4405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4409w4414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4409w4415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4419w4424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4419w4425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4429w4434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4429w4435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4439w4444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4439w4445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4449w4454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4449w4455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4459w4464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4459w4465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4469w4474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4469w4475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4479w4484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4479w4485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4209w4214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4209w4215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4489w4494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4489w4495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4499w4504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4499w4505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4509w4514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4509w4515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4519w4524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4519w4525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4529w4534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4529w4535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4539w4544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4539w4545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4549w4554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4549w4555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4559w4564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4559w4565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4569w4574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4569w4575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4579w4584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4579w4585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4219w4224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4219w4225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4589w4594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4589w4595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4599w4604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4599w4605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4609w4614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4609w4615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4619w4624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4619w4625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4629w4634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4629w4635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4639w4644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4639w4645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4649w4654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4649w4655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4659w4664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4659w4665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4669w4674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4669w4675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4679w4684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4679w4685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4229w4234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4229w4235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4689w4694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4689w4695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4699w4704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4699w4705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4709w4714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4709w4715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4719w4724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4719w4725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4729w4734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4729w4735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4739w4744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4739w4745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4749w4754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4749w4755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4759w4764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4759w4765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4769w4774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4769w4775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4779w4784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4779w4785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4239w4244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4239w4245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4789w4794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4789w4795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4799w4804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4799w4805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4809w4814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4809w4815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4819w4824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4819w4825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4829w4834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4829w4835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4839w4844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4839w4845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4849w4854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4849w4855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4859w4864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4859w4865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4869w4874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4869w4875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4879w4884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4879w4885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4249w4254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4249w4255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4889w4894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4889w4895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4899w4904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4899w4905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4909w4914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4909w4915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4919w4924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4919w4925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4929w4934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4929w4935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4939w4944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4939w4945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4949w4954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4949w4955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4959w4964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4959w4965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4969w4974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4969w4975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4979w4984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4979w4985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4259w4264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4259w4265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4989w4994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4989w4995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4999w5004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4999w5005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5009w5014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5009w5015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5019w5024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5019w5025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5029w5034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5029w5035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5039w5044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5039w5045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5049w5054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5049w5055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5059w5064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5059w5065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5069w5074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5069w5075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5079w5084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5079w5085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4269w4274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4269w4275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4279w4284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4279w4285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4184w4185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4124w4125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4118w4119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4112w4113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4106w4107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4100w4101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4094w4095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4088w4089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4082w4083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4076w4077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4070w4071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4178w4179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4064w4065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4058w4059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4052w4053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4046w4047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4040w4041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4034w4035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4028w4029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4022w4023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4016w4017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4010w4011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4172w4173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4004w4005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3998w3999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3992w3993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3986w3987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3980w3981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3974w3975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3968w3969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3962w3963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3956w3957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3950w3951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4166w4167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3944w3945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3938w3939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3932w3933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3926w3927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3920w3921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3914w3915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3908w3909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3902w3903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3896w3897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3890w3891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4160w4161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3884w3885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3878w3879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3872w3873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3866w3867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3860w3861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3854w3855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3848w3849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3842w3843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3836w3837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range3830w3831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4154w4155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4148w4149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4142w4143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4136w4137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lsb_prod_wo_range4130w4131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4181w4182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4121w4122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4115w4116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4109w4110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4103w4104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4097w4098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4091w4092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4085w4086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4079w4080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4073w4074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4067w4068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4175w4176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4061w4062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4055w4056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4049w4050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4043w4044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4037w4038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4031w4032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4025w4026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4019w4020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4013w4014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4007w4008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4169w4170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4001w4002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3995w3996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3989w3990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3983w3984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3977w3978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3971w3972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3965w3966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3959w3960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3953w3954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3947w3948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4163w4164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3941w3942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3935w3936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3929w3930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3923w3924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3917w3918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3911w3912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3905w3906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3899w3900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3893w3894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3887w3888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4157w4158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3881w3882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3875w3876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3869w3870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3863w3864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3857w3858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3851w3852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3845w3846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3839w3840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3833w3834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range3827w3828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4151w4152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4145w4146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4139w4140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4133w4134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_msb_prod_wo_range4127w4128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5094w5101w5102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5206w5212w5213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5217w5223w5224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5228w5234w5235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5239w5245w5246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5250w5256w5257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5261w5267w5268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5272w5278w5279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5283w5289w5290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5294w5300w5301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5305w5311w5312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5107w5113w5114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5316w5322w5323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5327w5333w5334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5338w5344w5345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5349w5355w5356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5360w5366w5367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5371w5377w5378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5382w5388w5389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5393w5399w5400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5404w5410w5411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5415w5421w5422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5118w5124w5125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5426w5432w5433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5437w5443w5444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5448w5454w5455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5459w5465w5466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5470w5476w5477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5481w5487w5488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5492w5498w5499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5503w5509w5510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5514w5520w5521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5525w5531w5532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5129w5135w5136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5536w5542w5543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5547w5553w5554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5558w5564w5565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5569w5575w5576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5580w5586w5587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5591w5597w5598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5602w5608w5609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5613w5619w5620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5624w5630w5631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5635w5641w5642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5140w5146w5147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5646w5652w5653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5657w5663w5664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5668w5674w5675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5679w5685w5686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5690w5696w5697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5701w5707w5708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5712w5718w5719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5723w5729w5730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5734w5740w5741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5745w5751w5752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5151w5157w5158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5756w5762w5763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5767w5773w5774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5778w5784w5785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5789w5795w5796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5800w5806w5807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5811w5817w5818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5822w5828w5829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5833w5839w5840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5844w5850w5851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5855w5861w5862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5162w5168w5169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5866w5872w5873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5877w5883w5884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5888w5894w5895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5899w5905w5906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5910w5916w5917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5921w5927w5928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5932w5938w5939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5943w5949w5950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5954w5960w5961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5965w5971w5972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5173w5179w5180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5976w5982w5983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5987w5993w5994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5998w6004w6005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6009w6015w6016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6020w6026w6027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6031w6037w6038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6042w6048w6049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6053w6059w6060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6064w6070w6071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6075w6081w6082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5184w5190w5191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5195w5201w5202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4187w4194w4195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4289w4295w4296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4299w4305w4306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4309w4315w4316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4319w4325w4326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4329w4335w4336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4339w4345w4346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4349w4355w4356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4359w4365w4366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4369w4375w4376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4379w4385w4386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4199w4205w4206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4389w4395w4396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4399w4405w4406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4409w4415w4416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4419w4425w4426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4429w4435w4436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4439w4445w4446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4449w4455w4456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4459w4465w4466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4469w4475w4476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4479w4485w4486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4209w4215w4216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4489w4495w4496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4499w4505w4506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4509w4515w4516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4519w4525w4526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4529w4535w4536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4539w4545w4546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4549w4555w4556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4559w4565w4566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4569w4575w4576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4579w4585w4586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4219w4225w4226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4589w4595w4596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4599w4605w4606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4609w4615w4616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4619w4625w4626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4629w4635w4636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4639w4645w4646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4649w4655w4656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4659w4665w4666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4669w4675w4676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4679w4685w4686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4229w4235w4236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4689w4695w4696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4699w4705w4706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4709w4715w4716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4719w4725w4726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4729w4735w4736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4739w4745w4746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4749w4755w4756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4759w4765w4766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4769w4775w4776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4779w4785w4786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4239w4245w4246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4789w4795w4796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4799w4805w4806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4809w4815w4816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4819w4825w4826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4829w4835w4836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4839w4845w4846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4849w4855w4856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4859w4865w4866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4869w4875w4876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4879w4885w4886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4249w4255w4256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4889w4895w4896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4899w4905w4906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4909w4915w4916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4919w4925w4926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4929w4935w4936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4939w4945w4946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4949w4955w4956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4959w4965w4966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4969w4975w4976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4979w4985w4986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4259w4265w4266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4989w4995w4996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4999w5005w5006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5009w5015w5016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5019w5025w5026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5029w5035w5036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5039w5045w5046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5049w5055w5056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5059w5065w5066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5069w5075w5076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5079w5085w5086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4269w4275w4276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4279w4285w4286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5094w5101w5102w5103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5206w5212w5213w5214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5217w5223w5224w5225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5228w5234w5235w5236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5239w5245w5246w5247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5250w5256w5257w5258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5261w5267w5268w5269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5272w5278w5279w5280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5283w5289w5290w5291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5294w5300w5301w5302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5305w5311w5312w5313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5107w5113w5114w5115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5316w5322w5323w5324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5327w5333w5334w5335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5338w5344w5345w5346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5349w5355w5356w5357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5360w5366w5367w5368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5371w5377w5378w5379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5382w5388w5389w5390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5393w5399w5400w5401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5404w5410w5411w5412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5415w5421w5422w5423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5118w5124w5125w5126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5426w5432w5433w5434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5437w5443w5444w5445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5448w5454w5455w5456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5459w5465w5466w5467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5470w5476w5477w5478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5481w5487w5488w5489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5492w5498w5499w5500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5503w5509w5510w5511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5514w5520w5521w5522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5525w5531w5532w5533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5129w5135w5136w5137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5536w5542w5543w5544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5547w5553w5554w5555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5558w5564w5565w5566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5569w5575w5576w5577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5580w5586w5587w5588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5591w5597w5598w5599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5602w5608w5609w5610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5613w5619w5620w5621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5624w5630w5631w5632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5635w5641w5642w5643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5140w5146w5147w5148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5646w5652w5653w5654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5657w5663w5664w5665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5668w5674w5675w5676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5679w5685w5686w5687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5690w5696w5697w5698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5701w5707w5708w5709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5712w5718w5719w5720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5723w5729w5730w5731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5734w5740w5741w5742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5745w5751w5752w5753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5151w5157w5158w5159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5756w5762w5763w5764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5767w5773w5774w5775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5778w5784w5785w5786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5789w5795w5796w5797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5800w5806w5807w5808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5811w5817w5818w5819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5822w5828w5829w5830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5833w5839w5840w5841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5844w5850w5851w5852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5855w5861w5862w5863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5162w5168w5169w5170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5866w5872w5873w5874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5877w5883w5884w5885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5888w5894w5895w5896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5899w5905w5906w5907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5910w5916w5917w5918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5921w5927w5928w5929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5932w5938w5939w5940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5943w5949w5950w5951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5954w5960w5961w5962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5965w5971w5972w5973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5173w5179w5180w5181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5976w5982w5983w5984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5987w5993w5994w5995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5998w6004w6005w6006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6009w6015w6016w6017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6020w6026w6027w6028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6031w6037w6038w6039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6042w6048w6049w6050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6053w6059w6060w6061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6064w6070w6071w6072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6075w6081w6082w6083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5184w5190w5191w5192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5195w5201w5202w5203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4187w4194w4195w4196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4289w4295w4296w4297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4299w4305w4306w4307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4309w4315w4316w4317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4319w4325w4326w4327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4329w4335w4336w4337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4339w4345w4346w4347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4349w4355w4356w4357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4359w4365w4366w4367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4369w4375w4376w4377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4379w4385w4386w4387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4199w4205w4206w4207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4389w4395w4396w4397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4399w4405w4406w4407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4409w4415w4416w4417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4419w4425w4426w4427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4429w4435w4436w4437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4439w4445w4446w4447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4449w4455w4456w4457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4459w4465w4466w4467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4469w4475w4476w4477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4479w4485w4486w4487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4209w4215w4216w4217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4489w4495w4496w4497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4499w4505w4506w4507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4509w4515w4516w4517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4519w4525w4526w4527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4529w4535w4536w4537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4539w4545w4546w4547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4549w4555w4556w4557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4559w4565w4566w4567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4569w4575w4576w4577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4579w4585w4586w4587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4219w4225w4226w4227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4589w4595w4596w4597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4599w4605w4606w4607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4609w4615w4616w4617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4619w4625w4626w4627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4629w4635w4636w4637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4639w4645w4646w4647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4649w4655w4656w4657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4659w4665w4666w4667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4669w4675w4676w4677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4679w4685w4686w4687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4229w4235w4236w4237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4689w4695w4696w4697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4699w4705w4706w4707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4709w4715w4716w4717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4719w4725w4726w4727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4729w4735w4736w4737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4739w4745w4746w4747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4749w4755w4756w4757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4759w4765w4766w4767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4769w4775w4776w4777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4779w4785w4786w4787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4239w4245w4246w4247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4789w4795w4796w4797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4799w4805w4806w4807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4809w4815w4816w4817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4819w4825w4826w4827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4829w4835w4836w4837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4839w4845w4846w4847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4849w4855w4856w4857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4859w4865w4866w4867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4869w4875w4876w4877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4879w4885w4886w4887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4249w4255w4256w4257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4889w4895w4896w4897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4899w4905w4906w4907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4909w4915w4916w4917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4919w4925w4926w4927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4929w4935w4936w4937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4939w4945w4946w4947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4949w4955w4956w4957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4959w4965w4966w4967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4969w4975w4976w4977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4979w4985w4986w4987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4259w4265w4266w4267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4989w4995w4996w4997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4999w5005w5006w5007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5009w5015w5016w5017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5019w5025w5026w5027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5029w5035w5036w5037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5039w5045w5046w5047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5049w5055w5056w5057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5059w5065w5066w5067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5069w5075w5076w5077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5079w5085w5086w5087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4269w4275w4276w4277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4279w4285w4286w4287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5094w5095w5096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5206w5207w5208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5217w5218w5219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5228w5229w5230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5239w5240w5241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5250w5251w5252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5261w5262w5263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5272w5273w5274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5283w5284w5285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5294w5295w5296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5305w5306w5307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5107w5108w5109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5316w5317w5318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5327w5328w5329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5338w5339w5340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5349w5350w5351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5360w5361w5362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5371w5372w5373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5382w5383w5384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5393w5394w5395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5404w5405w5406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5415w5416w5417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5118w5119w5120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5426w5427w5428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5437w5438w5439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5448w5449w5450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5459w5460w5461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5470w5471w5472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5481w5482w5483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5492w5493w5494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5503w5504w5505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5514w5515w5516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5525w5526w5527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5129w5130w5131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5536w5537w5538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5547w5548w5549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5558w5559w5560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5569w5570w5571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5580w5581w5582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5591w5592w5593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5602w5603w5604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5613w5614w5615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5624w5625w5626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5635w5636w5637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5140w5141w5142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5646w5647w5648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5657w5658w5659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5668w5669w5670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5679w5680w5681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5690w5691w5692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5701w5702w5703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5712w5713w5714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5723w5724w5725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5734w5735w5736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5745w5746w5747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5151w5152w5153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5756w5757w5758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5767w5768w5769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5778w5779w5780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5789w5790w5791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5800w5801w5802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5811w5812w5813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5822w5823w5824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5833w5834w5835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5844w5845w5846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5855w5856w5857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5162w5163w5164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5866w5867w5868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5877w5878w5879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5888w5889w5890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5899w5900w5901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5910w5911w5912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5921w5922w5923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5932w5933w5934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5943w5944w5945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5954w5955w5956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5965w5966w5967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5173w5174w5175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5976w5977w5978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5987w5988w5989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5998w5999w6000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6009w6010w6011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6020w6021w6022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6031w6032w6033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6042w6043w6044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6053w6054w6055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6064w6065w6066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range6075w6076w6077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5184w5185w5186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector1_range5195w5196w5197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4187w4188w4189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4289w4290w4291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4299w4300w4301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4309w4310w4311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4319w4320w4321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4329w4330w4331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4339w4340w4341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4349w4350w4351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4359w4360w4361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4369w4370w4371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4379w4380w4381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4199w4200w4201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4389w4390w4391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4399w4400w4401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4409w4410w4411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4419w4420w4421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4429w4430w4431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4439w4440w4441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4449w4450w4451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4459w4460w4461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4469w4470w4471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4479w4480w4481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4209w4210w4211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4489w4490w4491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4499w4500w4501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4509w4510w4511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4519w4520w4521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4529w4530w4531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4539w4540w4541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4549w4550w4551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4559w4560w4561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4569w4570w4571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4579w4580w4581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4219w4220w4221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4589w4590w4591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4599w4600w4601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4609w4610w4611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4619w4620w4621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4629w4630w4631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4639w4640w4641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4649w4650w4651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4659w4660w4661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4669w4670w4671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4679w4680w4681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4229w4230w4231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4689w4690w4691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4699w4700w4701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4709w4710w4711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4719w4720w4721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4729w4730w4731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4739w4740w4741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4749w4750w4751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4759w4760w4761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4769w4770w4771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4779w4780w4781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4239w4240w4241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4789w4790w4791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4799w4800w4801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4809w4810w4811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4819w4820w4821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4829w4830w4831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4839w4840w4841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4849w4850w4851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4859w4860w4861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4869w4870w4871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4879w4880w4881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4249w4250w4251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4889w4890w4891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4899w4900w4901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4909w4910w4911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4919w4920w4921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4929w4930w4931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4939w4940w4941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4949w4950w4951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4959w4960w4961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4969w4970w4971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4979w4980w4981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4259w4260w4261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4989w4990w4991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4999w5000w5001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5009w5010w5011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5019w5020w5021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5029w5030w5031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5039w5040w5041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5049w5050w5051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5059w5060w5061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5069w5070w5071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range5079w5080w5081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4269w4270w4271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_lg_w_vector2_range4279w4280w4281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5094w5095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5206w5207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5217w5218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5228w5229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5239w5240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5250w5251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5261w5262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5272w5273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5283w5284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5294w5295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5305w5306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5107w5108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5316w5317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5327w5328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5338w5339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5349w5350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5360w5361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5371w5372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5382w5383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5393w5394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5404w5405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5415w5416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5118w5119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5426w5427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5437w5438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5448w5449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5459w5460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5470w5471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5481w5482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5492w5493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5503w5504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5514w5515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5525w5526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5129w5130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5536w5537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5547w5548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5558w5559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5569w5570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5580w5581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5591w5592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5602w5603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5613w5614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5624w5625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5635w5636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5140w5141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5646w5647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5657w5658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5668w5669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5679w5680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5690w5691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5701w5702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5712w5713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5723w5724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5734w5735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5745w5746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5151w5152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5756w5757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5767w5768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5778w5779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5789w5790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5800w5801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5811w5812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5822w5823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5833w5834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5844w5845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5855w5856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5162w5163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5866w5867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5877w5878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5888w5889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5899w5900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5910w5911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5921w5922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5932w5933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5943w5944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5954w5955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5965w5966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5173w5174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5976w5977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5987w5988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5998w5999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6009w6010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6020w6021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6031w6032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6042w6043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6053w6054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6064w6065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range6075w6076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5184w5185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector1_range5195w5196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4187w4188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4289w4290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4299w4300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4309w4310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4319w4320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4329w4330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4339w4340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4349w4350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4359w4360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4369w4370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4379w4380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4199w4200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4389w4390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4399w4400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4409w4410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4419w4420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4429w4430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4439w4440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4449w4450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4459w4460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4469w4470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4479w4480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4209w4210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4489w4490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4499w4500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4509w4510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4519w4520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4529w4530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4539w4540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4549w4550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4559w4560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4569w4570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4579w4580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4219w4220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4589w4590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4599w4600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4609w4610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4619w4620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4629w4630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4639w4640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4649w4650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4659w4660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4669w4670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4679w4680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4229w4230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4689w4690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4699w4700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4709w4710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4719w4720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4729w4730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4739w4740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4749w4750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4759w4760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4769w4770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4779w4780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4239w4240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4789w4790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4799w4800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4809w4810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4819w4820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4829w4830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4839w4840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4849w4850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4859w4860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4869w4870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4879w4880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4249w4250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4889w4890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4899w4900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4909w4910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4919w4920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4929w4930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4939w4940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4949w4950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4959w4960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4969w4970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4979w4980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4259w4260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4989w4990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4999w5000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5009w5010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5019w5020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5029w5030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5039w5040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5049w5050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5059w5060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5069w5070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range5079w5080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4269w4270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lg_w_vector2_range4279w4280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  car_one :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_one_adj :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_two :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_two_adj :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_two_wo :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  lowest_bits_wi :	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  lowest_bits_wo :	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  lsb_prod_wi :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  lsb_prod_wo :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  mid_prod_wi :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  mid_prod_wo :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  msb_prod_out :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  msb_prod_wi :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  msb_prod_wo :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  neg_lsb :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  neg_msb :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  sum_one :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  sum_two :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  sum_two_wo :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  vector1 :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  vector2 :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  wire_a :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_b :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range6074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_car_one_adj_range5194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range3830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_lsb_prod_wo_range4130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range3827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_msb_prod_wo_range4127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range3708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_lsb_range4132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range3705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_neg_msb_range4129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range5082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_sum_one_range4282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range6075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector1_range5195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range5079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_prod_w_vector2_range4279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  ALTFP_EXa_altmult_opt_csa_ksf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(89 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(89 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(89 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_man_prod_w_lg_w_neg_msb_range4183w4192w(0) <= wire_man_prod_w_neg_msb_range4183w(0) AND wire_man_prod_w_neg_lsb_range4186w(0);
	wire_man_prod_w_lg_w_neg_msb_range4123w4293w(0) <= wire_man_prod_w_neg_msb_range4123w(0) AND wire_man_prod_w_neg_lsb_range4126w(0);
	wire_man_prod_w_lg_w_neg_msb_range4117w4303w(0) <= wire_man_prod_w_neg_msb_range4117w(0) AND wire_man_prod_w_neg_lsb_range4120w(0);
	wire_man_prod_w_lg_w_neg_msb_range4111w4313w(0) <= wire_man_prod_w_neg_msb_range4111w(0) AND wire_man_prod_w_neg_lsb_range4114w(0);
	wire_man_prod_w_lg_w_neg_msb_range4105w4323w(0) <= wire_man_prod_w_neg_msb_range4105w(0) AND wire_man_prod_w_neg_lsb_range4108w(0);
	wire_man_prod_w_lg_w_neg_msb_range4099w4333w(0) <= wire_man_prod_w_neg_msb_range4099w(0) AND wire_man_prod_w_neg_lsb_range4102w(0);
	wire_man_prod_w_lg_w_neg_msb_range4093w4343w(0) <= wire_man_prod_w_neg_msb_range4093w(0) AND wire_man_prod_w_neg_lsb_range4096w(0);
	wire_man_prod_w_lg_w_neg_msb_range4087w4353w(0) <= wire_man_prod_w_neg_msb_range4087w(0) AND wire_man_prod_w_neg_lsb_range4090w(0);
	wire_man_prod_w_lg_w_neg_msb_range4081w4363w(0) <= wire_man_prod_w_neg_msb_range4081w(0) AND wire_man_prod_w_neg_lsb_range4084w(0);
	wire_man_prod_w_lg_w_neg_msb_range4075w4373w(0) <= wire_man_prod_w_neg_msb_range4075w(0) AND wire_man_prod_w_neg_lsb_range4078w(0);
	wire_man_prod_w_lg_w_neg_msb_range4069w4383w(0) <= wire_man_prod_w_neg_msb_range4069w(0) AND wire_man_prod_w_neg_lsb_range4072w(0);
	wire_man_prod_w_lg_w_neg_msb_range4177w4203w(0) <= wire_man_prod_w_neg_msb_range4177w(0) AND wire_man_prod_w_neg_lsb_range4180w(0);
	wire_man_prod_w_lg_w_neg_msb_range4063w4393w(0) <= wire_man_prod_w_neg_msb_range4063w(0) AND wire_man_prod_w_neg_lsb_range4066w(0);
	wire_man_prod_w_lg_w_neg_msb_range4057w4403w(0) <= wire_man_prod_w_neg_msb_range4057w(0) AND wire_man_prod_w_neg_lsb_range4060w(0);
	wire_man_prod_w_lg_w_neg_msb_range4051w4413w(0) <= wire_man_prod_w_neg_msb_range4051w(0) AND wire_man_prod_w_neg_lsb_range4054w(0);
	wire_man_prod_w_lg_w_neg_msb_range4045w4423w(0) <= wire_man_prod_w_neg_msb_range4045w(0) AND wire_man_prod_w_neg_lsb_range4048w(0);
	wire_man_prod_w_lg_w_neg_msb_range4039w4433w(0) <= wire_man_prod_w_neg_msb_range4039w(0) AND wire_man_prod_w_neg_lsb_range4042w(0);
	wire_man_prod_w_lg_w_neg_msb_range4033w4443w(0) <= wire_man_prod_w_neg_msb_range4033w(0) AND wire_man_prod_w_neg_lsb_range4036w(0);
	wire_man_prod_w_lg_w_neg_msb_range4027w4453w(0) <= wire_man_prod_w_neg_msb_range4027w(0) AND wire_man_prod_w_neg_lsb_range4030w(0);
	wire_man_prod_w_lg_w_neg_msb_range4021w4463w(0) <= wire_man_prod_w_neg_msb_range4021w(0) AND wire_man_prod_w_neg_lsb_range4024w(0);
	wire_man_prod_w_lg_w_neg_msb_range4015w4473w(0) <= wire_man_prod_w_neg_msb_range4015w(0) AND wire_man_prod_w_neg_lsb_range4018w(0);
	wire_man_prod_w_lg_w_neg_msb_range4009w4483w(0) <= wire_man_prod_w_neg_msb_range4009w(0) AND wire_man_prod_w_neg_lsb_range4012w(0);
	wire_man_prod_w_lg_w_neg_msb_range4171w4213w(0) <= wire_man_prod_w_neg_msb_range4171w(0) AND wire_man_prod_w_neg_lsb_range4174w(0);
	wire_man_prod_w_lg_w_neg_msb_range4003w4493w(0) <= wire_man_prod_w_neg_msb_range4003w(0) AND wire_man_prod_w_neg_lsb_range4006w(0);
	wire_man_prod_w_lg_w_neg_msb_range3997w4503w(0) <= wire_man_prod_w_neg_msb_range3997w(0) AND wire_man_prod_w_neg_lsb_range4000w(0);
	wire_man_prod_w_lg_w_neg_msb_range3991w4513w(0) <= wire_man_prod_w_neg_msb_range3991w(0) AND wire_man_prod_w_neg_lsb_range3994w(0);
	wire_man_prod_w_lg_w_neg_msb_range3985w4523w(0) <= wire_man_prod_w_neg_msb_range3985w(0) AND wire_man_prod_w_neg_lsb_range3988w(0);
	wire_man_prod_w_lg_w_neg_msb_range3979w4533w(0) <= wire_man_prod_w_neg_msb_range3979w(0) AND wire_man_prod_w_neg_lsb_range3982w(0);
	wire_man_prod_w_lg_w_neg_msb_range3973w4543w(0) <= wire_man_prod_w_neg_msb_range3973w(0) AND wire_man_prod_w_neg_lsb_range3976w(0);
	wire_man_prod_w_lg_w_neg_msb_range3967w4553w(0) <= wire_man_prod_w_neg_msb_range3967w(0) AND wire_man_prod_w_neg_lsb_range3970w(0);
	wire_man_prod_w_lg_w_neg_msb_range3961w4563w(0) <= wire_man_prod_w_neg_msb_range3961w(0) AND wire_man_prod_w_neg_lsb_range3964w(0);
	wire_man_prod_w_lg_w_neg_msb_range3955w4573w(0) <= wire_man_prod_w_neg_msb_range3955w(0) AND wire_man_prod_w_neg_lsb_range3958w(0);
	wire_man_prod_w_lg_w_neg_msb_range3949w4583w(0) <= wire_man_prod_w_neg_msb_range3949w(0) AND wire_man_prod_w_neg_lsb_range3952w(0);
	wire_man_prod_w_lg_w_neg_msb_range4165w4223w(0) <= wire_man_prod_w_neg_msb_range4165w(0) AND wire_man_prod_w_neg_lsb_range4168w(0);
	wire_man_prod_w_lg_w_neg_msb_range3943w4593w(0) <= wire_man_prod_w_neg_msb_range3943w(0) AND wire_man_prod_w_neg_lsb_range3946w(0);
	wire_man_prod_w_lg_w_neg_msb_range3937w4603w(0) <= wire_man_prod_w_neg_msb_range3937w(0) AND wire_man_prod_w_neg_lsb_range3940w(0);
	wire_man_prod_w_lg_w_neg_msb_range3931w4613w(0) <= wire_man_prod_w_neg_msb_range3931w(0) AND wire_man_prod_w_neg_lsb_range3934w(0);
	wire_man_prod_w_lg_w_neg_msb_range3925w4623w(0) <= wire_man_prod_w_neg_msb_range3925w(0) AND wire_man_prod_w_neg_lsb_range3928w(0);
	wire_man_prod_w_lg_w_neg_msb_range3919w4633w(0) <= wire_man_prod_w_neg_msb_range3919w(0) AND wire_man_prod_w_neg_lsb_range3922w(0);
	wire_man_prod_w_lg_w_neg_msb_range3913w4643w(0) <= wire_man_prod_w_neg_msb_range3913w(0) AND wire_man_prod_w_neg_lsb_range3916w(0);
	wire_man_prod_w_lg_w_neg_msb_range3907w4653w(0) <= wire_man_prod_w_neg_msb_range3907w(0) AND wire_man_prod_w_neg_lsb_range3910w(0);
	wire_man_prod_w_lg_w_neg_msb_range3901w4663w(0) <= wire_man_prod_w_neg_msb_range3901w(0) AND wire_man_prod_w_neg_lsb_range3904w(0);
	wire_man_prod_w_lg_w_neg_msb_range3895w4673w(0) <= wire_man_prod_w_neg_msb_range3895w(0) AND wire_man_prod_w_neg_lsb_range3898w(0);
	wire_man_prod_w_lg_w_neg_msb_range3889w4683w(0) <= wire_man_prod_w_neg_msb_range3889w(0) AND wire_man_prod_w_neg_lsb_range3892w(0);
	wire_man_prod_w_lg_w_neg_msb_range4159w4233w(0) <= wire_man_prod_w_neg_msb_range4159w(0) AND wire_man_prod_w_neg_lsb_range4162w(0);
	wire_man_prod_w_lg_w_neg_msb_range3883w4693w(0) <= wire_man_prod_w_neg_msb_range3883w(0) AND wire_man_prod_w_neg_lsb_range3886w(0);
	wire_man_prod_w_lg_w_neg_msb_range3877w4703w(0) <= wire_man_prod_w_neg_msb_range3877w(0) AND wire_man_prod_w_neg_lsb_range3880w(0);
	wire_man_prod_w_lg_w_neg_msb_range3871w4713w(0) <= wire_man_prod_w_neg_msb_range3871w(0) AND wire_man_prod_w_neg_lsb_range3874w(0);
	wire_man_prod_w_lg_w_neg_msb_range3865w4723w(0) <= wire_man_prod_w_neg_msb_range3865w(0) AND wire_man_prod_w_neg_lsb_range3868w(0);
	wire_man_prod_w_lg_w_neg_msb_range3859w4733w(0) <= wire_man_prod_w_neg_msb_range3859w(0) AND wire_man_prod_w_neg_lsb_range3862w(0);
	wire_man_prod_w_lg_w_neg_msb_range3853w4743w(0) <= wire_man_prod_w_neg_msb_range3853w(0) AND wire_man_prod_w_neg_lsb_range3856w(0);
	wire_man_prod_w_lg_w_neg_msb_range3847w4753w(0) <= wire_man_prod_w_neg_msb_range3847w(0) AND wire_man_prod_w_neg_lsb_range3850w(0);
	wire_man_prod_w_lg_w_neg_msb_range3841w4763w(0) <= wire_man_prod_w_neg_msb_range3841w(0) AND wire_man_prod_w_neg_lsb_range3844w(0);
	wire_man_prod_w_lg_w_neg_msb_range3835w4773w(0) <= wire_man_prod_w_neg_msb_range3835w(0) AND wire_man_prod_w_neg_lsb_range3838w(0);
	wire_man_prod_w_lg_w_neg_msb_range3829w4783w(0) <= wire_man_prod_w_neg_msb_range3829w(0) AND wire_man_prod_w_neg_lsb_range3832w(0);
	wire_man_prod_w_lg_w_neg_msb_range4153w4243w(0) <= wire_man_prod_w_neg_msb_range4153w(0) AND wire_man_prod_w_neg_lsb_range4156w(0);
	wire_man_prod_w_lg_w_neg_msb_range3823w4793w(0) <= wire_man_prod_w_neg_msb_range3823w(0) AND wire_man_prod_w_neg_lsb_range3825w(0);
	wire_man_prod_w_lg_w_neg_msb_range3819w4803w(0) <= wire_man_prod_w_neg_msb_range3819w(0) AND wire_man_prod_w_neg_lsb_range3821w(0);
	wire_man_prod_w_lg_w_neg_msb_range3815w4813w(0) <= wire_man_prod_w_neg_msb_range3815w(0) AND wire_man_prod_w_neg_lsb_range3817w(0);
	wire_man_prod_w_lg_w_neg_msb_range3811w4823w(0) <= wire_man_prod_w_neg_msb_range3811w(0) AND wire_man_prod_w_neg_lsb_range3813w(0);
	wire_man_prod_w_lg_w_neg_msb_range3807w4833w(0) <= wire_man_prod_w_neg_msb_range3807w(0) AND wire_man_prod_w_neg_lsb_range3809w(0);
	wire_man_prod_w_lg_w_neg_msb_range3803w4843w(0) <= wire_man_prod_w_neg_msb_range3803w(0) AND wire_man_prod_w_neg_lsb_range3805w(0);
	wire_man_prod_w_lg_w_neg_msb_range3799w4853w(0) <= wire_man_prod_w_neg_msb_range3799w(0) AND wire_man_prod_w_neg_lsb_range3801w(0);
	wire_man_prod_w_lg_w_neg_msb_range3795w4863w(0) <= wire_man_prod_w_neg_msb_range3795w(0) AND wire_man_prod_w_neg_lsb_range3797w(0);
	wire_man_prod_w_lg_w_neg_msb_range3791w4873w(0) <= wire_man_prod_w_neg_msb_range3791w(0) AND wire_man_prod_w_neg_lsb_range3793w(0);
	wire_man_prod_w_lg_w_neg_msb_range3787w4883w(0) <= wire_man_prod_w_neg_msb_range3787w(0) AND wire_man_prod_w_neg_lsb_range3789w(0);
	wire_man_prod_w_lg_w_neg_msb_range4147w4253w(0) <= wire_man_prod_w_neg_msb_range4147w(0) AND wire_man_prod_w_neg_lsb_range4150w(0);
	wire_man_prod_w_lg_w_neg_msb_range3783w4893w(0) <= wire_man_prod_w_neg_msb_range3783w(0) AND wire_man_prod_w_neg_lsb_range3785w(0);
	wire_man_prod_w_lg_w_neg_msb_range3779w4903w(0) <= wire_man_prod_w_neg_msb_range3779w(0) AND wire_man_prod_w_neg_lsb_range3781w(0);
	wire_man_prod_w_lg_w_neg_msb_range3775w4913w(0) <= wire_man_prod_w_neg_msb_range3775w(0) AND wire_man_prod_w_neg_lsb_range3777w(0);
	wire_man_prod_w_lg_w_neg_msb_range3771w4923w(0) <= wire_man_prod_w_neg_msb_range3771w(0) AND wire_man_prod_w_neg_lsb_range3773w(0);
	wire_man_prod_w_lg_w_neg_msb_range3767w4933w(0) <= wire_man_prod_w_neg_msb_range3767w(0) AND wire_man_prod_w_neg_lsb_range3769w(0);
	wire_man_prod_w_lg_w_neg_msb_range3763w4943w(0) <= wire_man_prod_w_neg_msb_range3763w(0) AND wire_man_prod_w_neg_lsb_range3765w(0);
	wire_man_prod_w_lg_w_neg_msb_range3759w4953w(0) <= wire_man_prod_w_neg_msb_range3759w(0) AND wire_man_prod_w_neg_lsb_range3761w(0);
	wire_man_prod_w_lg_w_neg_msb_range3755w4963w(0) <= wire_man_prod_w_neg_msb_range3755w(0) AND wire_man_prod_w_neg_lsb_range3757w(0);
	wire_man_prod_w_lg_w_neg_msb_range3751w4973w(0) <= wire_man_prod_w_neg_msb_range3751w(0) AND wire_man_prod_w_neg_lsb_range3753w(0);
	wire_man_prod_w_lg_w_neg_msb_range3747w4983w(0) <= wire_man_prod_w_neg_msb_range3747w(0) AND wire_man_prod_w_neg_lsb_range3749w(0);
	wire_man_prod_w_lg_w_neg_msb_range4141w4263w(0) <= wire_man_prod_w_neg_msb_range4141w(0) AND wire_man_prod_w_neg_lsb_range4144w(0);
	wire_man_prod_w_lg_w_neg_msb_range3743w4993w(0) <= wire_man_prod_w_neg_msb_range3743w(0) AND wire_man_prod_w_neg_lsb_range3745w(0);
	wire_man_prod_w_lg_w_neg_msb_range3739w5003w(0) <= wire_man_prod_w_neg_msb_range3739w(0) AND wire_man_prod_w_neg_lsb_range3741w(0);
	wire_man_prod_w_lg_w_neg_msb_range3735w5013w(0) <= wire_man_prod_w_neg_msb_range3735w(0) AND wire_man_prod_w_neg_lsb_range3737w(0);
	wire_man_prod_w_lg_w_neg_msb_range3731w5023w(0) <= wire_man_prod_w_neg_msb_range3731w(0) AND wire_man_prod_w_neg_lsb_range3733w(0);
	wire_man_prod_w_lg_w_neg_msb_range3727w5033w(0) <= wire_man_prod_w_neg_msb_range3727w(0) AND wire_man_prod_w_neg_lsb_range3729w(0);
	wire_man_prod_w_lg_w_neg_msb_range3723w5043w(0) <= wire_man_prod_w_neg_msb_range3723w(0) AND wire_man_prod_w_neg_lsb_range3725w(0);
	wire_man_prod_w_lg_w_neg_msb_range3719w5053w(0) <= wire_man_prod_w_neg_msb_range3719w(0) AND wire_man_prod_w_neg_lsb_range3721w(0);
	wire_man_prod_w_lg_w_neg_msb_range3715w5063w(0) <= wire_man_prod_w_neg_msb_range3715w(0) AND wire_man_prod_w_neg_lsb_range3717w(0);
	wire_man_prod_w_lg_w_neg_msb_range3711w5073w(0) <= wire_man_prod_w_neg_msb_range3711w(0) AND wire_man_prod_w_neg_lsb_range3713w(0);
	wire_man_prod_w_lg_w_neg_msb_range3705w5083w(0) <= wire_man_prod_w_neg_msb_range3705w(0) AND wire_man_prod_w_neg_lsb_range3708w(0);
	wire_man_prod_w_lg_w_neg_msb_range4135w4273w(0) <= wire_man_prod_w_neg_msb_range4135w(0) AND wire_man_prod_w_neg_lsb_range4138w(0);
	wire_man_prod_w_lg_w_neg_msb_range4129w4283w(0) <= wire_man_prod_w_neg_msb_range4129w(0) AND wire_man_prod_w_neg_lsb_range4132w(0);
	wire_man_prod_w_lg_w_sum_one_range4190w5099w(0) <= wire_man_prod_w_sum_one_range4190w(0) AND wire_man_prod_w_car_one_adj_range5092w(0);
	wire_man_prod_w_lg_w_sum_one_range4292w5210w(0) <= wire_man_prod_w_sum_one_range4292w(0) AND wire_man_prod_w_car_one_adj_range5205w(0);
	wire_man_prod_w_lg_w_sum_one_range4302w5221w(0) <= wire_man_prod_w_sum_one_range4302w(0) AND wire_man_prod_w_car_one_adj_range5216w(0);
	wire_man_prod_w_lg_w_sum_one_range4312w5232w(0) <= wire_man_prod_w_sum_one_range4312w(0) AND wire_man_prod_w_car_one_adj_range5227w(0);
	wire_man_prod_w_lg_w_sum_one_range4322w5243w(0) <= wire_man_prod_w_sum_one_range4322w(0) AND wire_man_prod_w_car_one_adj_range5238w(0);
	wire_man_prod_w_lg_w_sum_one_range4332w5254w(0) <= wire_man_prod_w_sum_one_range4332w(0) AND wire_man_prod_w_car_one_adj_range5249w(0);
	wire_man_prod_w_lg_w_sum_one_range4342w5265w(0) <= wire_man_prod_w_sum_one_range4342w(0) AND wire_man_prod_w_car_one_adj_range5260w(0);
	wire_man_prod_w_lg_w_sum_one_range4352w5276w(0) <= wire_man_prod_w_sum_one_range4352w(0) AND wire_man_prod_w_car_one_adj_range5271w(0);
	wire_man_prod_w_lg_w_sum_one_range4362w5287w(0) <= wire_man_prod_w_sum_one_range4362w(0) AND wire_man_prod_w_car_one_adj_range5282w(0);
	wire_man_prod_w_lg_w_sum_one_range4372w5298w(0) <= wire_man_prod_w_sum_one_range4372w(0) AND wire_man_prod_w_car_one_adj_range5293w(0);
	wire_man_prod_w_lg_w_sum_one_range4382w5309w(0) <= wire_man_prod_w_sum_one_range4382w(0) AND wire_man_prod_w_car_one_adj_range5304w(0);
	wire_man_prod_w_lg_w_sum_one_range4202w5111w(0) <= wire_man_prod_w_sum_one_range4202w(0) AND wire_man_prod_w_car_one_adj_range5106w(0);
	wire_man_prod_w_lg_w_sum_one_range4392w5320w(0) <= wire_man_prod_w_sum_one_range4392w(0) AND wire_man_prod_w_car_one_adj_range5315w(0);
	wire_man_prod_w_lg_w_sum_one_range4402w5331w(0) <= wire_man_prod_w_sum_one_range4402w(0) AND wire_man_prod_w_car_one_adj_range5326w(0);
	wire_man_prod_w_lg_w_sum_one_range4412w5342w(0) <= wire_man_prod_w_sum_one_range4412w(0) AND wire_man_prod_w_car_one_adj_range5337w(0);
	wire_man_prod_w_lg_w_sum_one_range4422w5353w(0) <= wire_man_prod_w_sum_one_range4422w(0) AND wire_man_prod_w_car_one_adj_range5348w(0);
	wire_man_prod_w_lg_w_sum_one_range4432w5364w(0) <= wire_man_prod_w_sum_one_range4432w(0) AND wire_man_prod_w_car_one_adj_range5359w(0);
	wire_man_prod_w_lg_w_sum_one_range4442w5375w(0) <= wire_man_prod_w_sum_one_range4442w(0) AND wire_man_prod_w_car_one_adj_range5370w(0);
	wire_man_prod_w_lg_w_sum_one_range4452w5386w(0) <= wire_man_prod_w_sum_one_range4452w(0) AND wire_man_prod_w_car_one_adj_range5381w(0);
	wire_man_prod_w_lg_w_sum_one_range4462w5397w(0) <= wire_man_prod_w_sum_one_range4462w(0) AND wire_man_prod_w_car_one_adj_range5392w(0);
	wire_man_prod_w_lg_w_sum_one_range4472w5408w(0) <= wire_man_prod_w_sum_one_range4472w(0) AND wire_man_prod_w_car_one_adj_range5403w(0);
	wire_man_prod_w_lg_w_sum_one_range4482w5419w(0) <= wire_man_prod_w_sum_one_range4482w(0) AND wire_man_prod_w_car_one_adj_range5414w(0);
	wire_man_prod_w_lg_w_sum_one_range4212w5122w(0) <= wire_man_prod_w_sum_one_range4212w(0) AND wire_man_prod_w_car_one_adj_range5117w(0);
	wire_man_prod_w_lg_w_sum_one_range4492w5430w(0) <= wire_man_prod_w_sum_one_range4492w(0) AND wire_man_prod_w_car_one_adj_range5425w(0);
	wire_man_prod_w_lg_w_sum_one_range4502w5441w(0) <= wire_man_prod_w_sum_one_range4502w(0) AND wire_man_prod_w_car_one_adj_range5436w(0);
	wire_man_prod_w_lg_w_sum_one_range4512w5452w(0) <= wire_man_prod_w_sum_one_range4512w(0) AND wire_man_prod_w_car_one_adj_range5447w(0);
	wire_man_prod_w_lg_w_sum_one_range4522w5463w(0) <= wire_man_prod_w_sum_one_range4522w(0) AND wire_man_prod_w_car_one_adj_range5458w(0);
	wire_man_prod_w_lg_w_sum_one_range4532w5474w(0) <= wire_man_prod_w_sum_one_range4532w(0) AND wire_man_prod_w_car_one_adj_range5469w(0);
	wire_man_prod_w_lg_w_sum_one_range4542w5485w(0) <= wire_man_prod_w_sum_one_range4542w(0) AND wire_man_prod_w_car_one_adj_range5480w(0);
	wire_man_prod_w_lg_w_sum_one_range4552w5496w(0) <= wire_man_prod_w_sum_one_range4552w(0) AND wire_man_prod_w_car_one_adj_range5491w(0);
	wire_man_prod_w_lg_w_sum_one_range4562w5507w(0) <= wire_man_prod_w_sum_one_range4562w(0) AND wire_man_prod_w_car_one_adj_range5502w(0);
	wire_man_prod_w_lg_w_sum_one_range4572w5518w(0) <= wire_man_prod_w_sum_one_range4572w(0) AND wire_man_prod_w_car_one_adj_range5513w(0);
	wire_man_prod_w_lg_w_sum_one_range4582w5529w(0) <= wire_man_prod_w_sum_one_range4582w(0) AND wire_man_prod_w_car_one_adj_range5524w(0);
	wire_man_prod_w_lg_w_sum_one_range4222w5133w(0) <= wire_man_prod_w_sum_one_range4222w(0) AND wire_man_prod_w_car_one_adj_range5128w(0);
	wire_man_prod_w_lg_w_sum_one_range4592w5540w(0) <= wire_man_prod_w_sum_one_range4592w(0) AND wire_man_prod_w_car_one_adj_range5535w(0);
	wire_man_prod_w_lg_w_sum_one_range4602w5551w(0) <= wire_man_prod_w_sum_one_range4602w(0) AND wire_man_prod_w_car_one_adj_range5546w(0);
	wire_man_prod_w_lg_w_sum_one_range4612w5562w(0) <= wire_man_prod_w_sum_one_range4612w(0) AND wire_man_prod_w_car_one_adj_range5557w(0);
	wire_man_prod_w_lg_w_sum_one_range4622w5573w(0) <= wire_man_prod_w_sum_one_range4622w(0) AND wire_man_prod_w_car_one_adj_range5568w(0);
	wire_man_prod_w_lg_w_sum_one_range4632w5584w(0) <= wire_man_prod_w_sum_one_range4632w(0) AND wire_man_prod_w_car_one_adj_range5579w(0);
	wire_man_prod_w_lg_w_sum_one_range4642w5595w(0) <= wire_man_prod_w_sum_one_range4642w(0) AND wire_man_prod_w_car_one_adj_range5590w(0);
	wire_man_prod_w_lg_w_sum_one_range4652w5606w(0) <= wire_man_prod_w_sum_one_range4652w(0) AND wire_man_prod_w_car_one_adj_range5601w(0);
	wire_man_prod_w_lg_w_sum_one_range4662w5617w(0) <= wire_man_prod_w_sum_one_range4662w(0) AND wire_man_prod_w_car_one_adj_range5612w(0);
	wire_man_prod_w_lg_w_sum_one_range4672w5628w(0) <= wire_man_prod_w_sum_one_range4672w(0) AND wire_man_prod_w_car_one_adj_range5623w(0);
	wire_man_prod_w_lg_w_sum_one_range4682w5639w(0) <= wire_man_prod_w_sum_one_range4682w(0) AND wire_man_prod_w_car_one_adj_range5634w(0);
	wire_man_prod_w_lg_w_sum_one_range4232w5144w(0) <= wire_man_prod_w_sum_one_range4232w(0) AND wire_man_prod_w_car_one_adj_range5139w(0);
	wire_man_prod_w_lg_w_sum_one_range4692w5650w(0) <= wire_man_prod_w_sum_one_range4692w(0) AND wire_man_prod_w_car_one_adj_range5645w(0);
	wire_man_prod_w_lg_w_sum_one_range4702w5661w(0) <= wire_man_prod_w_sum_one_range4702w(0) AND wire_man_prod_w_car_one_adj_range5656w(0);
	wire_man_prod_w_lg_w_sum_one_range4712w5672w(0) <= wire_man_prod_w_sum_one_range4712w(0) AND wire_man_prod_w_car_one_adj_range5667w(0);
	wire_man_prod_w_lg_w_sum_one_range4722w5683w(0) <= wire_man_prod_w_sum_one_range4722w(0) AND wire_man_prod_w_car_one_adj_range5678w(0);
	wire_man_prod_w_lg_w_sum_one_range4732w5694w(0) <= wire_man_prod_w_sum_one_range4732w(0) AND wire_man_prod_w_car_one_adj_range5689w(0);
	wire_man_prod_w_lg_w_sum_one_range4742w5705w(0) <= wire_man_prod_w_sum_one_range4742w(0) AND wire_man_prod_w_car_one_adj_range5700w(0);
	wire_man_prod_w_lg_w_sum_one_range4752w5716w(0) <= wire_man_prod_w_sum_one_range4752w(0) AND wire_man_prod_w_car_one_adj_range5711w(0);
	wire_man_prod_w_lg_w_sum_one_range4762w5727w(0) <= wire_man_prod_w_sum_one_range4762w(0) AND wire_man_prod_w_car_one_adj_range5722w(0);
	wire_man_prod_w_lg_w_sum_one_range4772w5738w(0) <= wire_man_prod_w_sum_one_range4772w(0) AND wire_man_prod_w_car_one_adj_range5733w(0);
	wire_man_prod_w_lg_w_sum_one_range4782w5749w(0) <= wire_man_prod_w_sum_one_range4782w(0) AND wire_man_prod_w_car_one_adj_range5744w(0);
	wire_man_prod_w_lg_w_sum_one_range4242w5155w(0) <= wire_man_prod_w_sum_one_range4242w(0) AND wire_man_prod_w_car_one_adj_range5150w(0);
	wire_man_prod_w_lg_w_sum_one_range4792w5760w(0) <= wire_man_prod_w_sum_one_range4792w(0) AND wire_man_prod_w_car_one_adj_range5755w(0);
	wire_man_prod_w_lg_w_sum_one_range4802w5771w(0) <= wire_man_prod_w_sum_one_range4802w(0) AND wire_man_prod_w_car_one_adj_range5766w(0);
	wire_man_prod_w_lg_w_sum_one_range4812w5782w(0) <= wire_man_prod_w_sum_one_range4812w(0) AND wire_man_prod_w_car_one_adj_range5777w(0);
	wire_man_prod_w_lg_w_sum_one_range4822w5793w(0) <= wire_man_prod_w_sum_one_range4822w(0) AND wire_man_prod_w_car_one_adj_range5788w(0);
	wire_man_prod_w_lg_w_sum_one_range4832w5804w(0) <= wire_man_prod_w_sum_one_range4832w(0) AND wire_man_prod_w_car_one_adj_range5799w(0);
	wire_man_prod_w_lg_w_sum_one_range4842w5815w(0) <= wire_man_prod_w_sum_one_range4842w(0) AND wire_man_prod_w_car_one_adj_range5810w(0);
	wire_man_prod_w_lg_w_sum_one_range4852w5826w(0) <= wire_man_prod_w_sum_one_range4852w(0) AND wire_man_prod_w_car_one_adj_range5821w(0);
	wire_man_prod_w_lg_w_sum_one_range4862w5837w(0) <= wire_man_prod_w_sum_one_range4862w(0) AND wire_man_prod_w_car_one_adj_range5832w(0);
	wire_man_prod_w_lg_w_sum_one_range4872w5848w(0) <= wire_man_prod_w_sum_one_range4872w(0) AND wire_man_prod_w_car_one_adj_range5843w(0);
	wire_man_prod_w_lg_w_sum_one_range4882w5859w(0) <= wire_man_prod_w_sum_one_range4882w(0) AND wire_man_prod_w_car_one_adj_range5854w(0);
	wire_man_prod_w_lg_w_sum_one_range4252w5166w(0) <= wire_man_prod_w_sum_one_range4252w(0) AND wire_man_prod_w_car_one_adj_range5161w(0);
	wire_man_prod_w_lg_w_sum_one_range4892w5870w(0) <= wire_man_prod_w_sum_one_range4892w(0) AND wire_man_prod_w_car_one_adj_range5865w(0);
	wire_man_prod_w_lg_w_sum_one_range4902w5881w(0) <= wire_man_prod_w_sum_one_range4902w(0) AND wire_man_prod_w_car_one_adj_range5876w(0);
	wire_man_prod_w_lg_w_sum_one_range4912w5892w(0) <= wire_man_prod_w_sum_one_range4912w(0) AND wire_man_prod_w_car_one_adj_range5887w(0);
	wire_man_prod_w_lg_w_sum_one_range4922w5903w(0) <= wire_man_prod_w_sum_one_range4922w(0) AND wire_man_prod_w_car_one_adj_range5898w(0);
	wire_man_prod_w_lg_w_sum_one_range4932w5914w(0) <= wire_man_prod_w_sum_one_range4932w(0) AND wire_man_prod_w_car_one_adj_range5909w(0);
	wire_man_prod_w_lg_w_sum_one_range4942w5925w(0) <= wire_man_prod_w_sum_one_range4942w(0) AND wire_man_prod_w_car_one_adj_range5920w(0);
	wire_man_prod_w_lg_w_sum_one_range4952w5936w(0) <= wire_man_prod_w_sum_one_range4952w(0) AND wire_man_prod_w_car_one_adj_range5931w(0);
	wire_man_prod_w_lg_w_sum_one_range4962w5947w(0) <= wire_man_prod_w_sum_one_range4962w(0) AND wire_man_prod_w_car_one_adj_range5942w(0);
	wire_man_prod_w_lg_w_sum_one_range4972w5958w(0) <= wire_man_prod_w_sum_one_range4972w(0) AND wire_man_prod_w_car_one_adj_range5953w(0);
	wire_man_prod_w_lg_w_sum_one_range4982w5969w(0) <= wire_man_prod_w_sum_one_range4982w(0) AND wire_man_prod_w_car_one_adj_range5964w(0);
	wire_man_prod_w_lg_w_sum_one_range4262w5177w(0) <= wire_man_prod_w_sum_one_range4262w(0) AND wire_man_prod_w_car_one_adj_range5172w(0);
	wire_man_prod_w_lg_w_sum_one_range4992w5980w(0) <= wire_man_prod_w_sum_one_range4992w(0) AND wire_man_prod_w_car_one_adj_range5975w(0);
	wire_man_prod_w_lg_w_sum_one_range5002w5991w(0) <= wire_man_prod_w_sum_one_range5002w(0) AND wire_man_prod_w_car_one_adj_range5986w(0);
	wire_man_prod_w_lg_w_sum_one_range5012w6002w(0) <= wire_man_prod_w_sum_one_range5012w(0) AND wire_man_prod_w_car_one_adj_range5997w(0);
	wire_man_prod_w_lg_w_sum_one_range5022w6013w(0) <= wire_man_prod_w_sum_one_range5022w(0) AND wire_man_prod_w_car_one_adj_range6008w(0);
	wire_man_prod_w_lg_w_sum_one_range5032w6024w(0) <= wire_man_prod_w_sum_one_range5032w(0) AND wire_man_prod_w_car_one_adj_range6019w(0);
	wire_man_prod_w_lg_w_sum_one_range5042w6035w(0) <= wire_man_prod_w_sum_one_range5042w(0) AND wire_man_prod_w_car_one_adj_range6030w(0);
	wire_man_prod_w_lg_w_sum_one_range5052w6046w(0) <= wire_man_prod_w_sum_one_range5052w(0) AND wire_man_prod_w_car_one_adj_range6041w(0);
	wire_man_prod_w_lg_w_sum_one_range5062w6057w(0) <= wire_man_prod_w_sum_one_range5062w(0) AND wire_man_prod_w_car_one_adj_range6052w(0);
	wire_man_prod_w_lg_w_sum_one_range5072w6068w(0) <= wire_man_prod_w_sum_one_range5072w(0) AND wire_man_prod_w_car_one_adj_range6063w(0);
	wire_man_prod_w_lg_w_sum_one_range5082w6079w(0) <= wire_man_prod_w_sum_one_range5082w(0) AND wire_man_prod_w_car_one_adj_range6074w(0);
	wire_man_prod_w_lg_w_sum_one_range4272w5188w(0) <= wire_man_prod_w_sum_one_range4272w(0) AND wire_man_prod_w_car_one_adj_range5183w(0);
	wire_man_prod_w_lg_w_sum_one_range4282w5199w(0) <= wire_man_prod_w_sum_one_range4282w(0) AND wire_man_prod_w_car_one_adj_range5194w(0);
	wire_man_prod_w_lg_w_vector1_range5094w5100w(0) <= wire_man_prod_w_vector1_range5094w(0) AND wire_man_prod_w_car_one_adj_range5092w(0);
	wire_man_prod_w_lg_w_vector1_range5094w5101w(0) <= wire_man_prod_w_vector1_range5094w(0) AND wire_man_prod_w_sum_one_range4190w(0);
	wire_man_prod_w_lg_w_vector1_range5206w5211w(0) <= wire_man_prod_w_vector1_range5206w(0) AND wire_man_prod_w_car_one_adj_range5205w(0);
	wire_man_prod_w_lg_w_vector1_range5206w5212w(0) <= wire_man_prod_w_vector1_range5206w(0) AND wire_man_prod_w_sum_one_range4292w(0);
	wire_man_prod_w_lg_w_vector1_range5217w5222w(0) <= wire_man_prod_w_vector1_range5217w(0) AND wire_man_prod_w_car_one_adj_range5216w(0);
	wire_man_prod_w_lg_w_vector1_range5217w5223w(0) <= wire_man_prod_w_vector1_range5217w(0) AND wire_man_prod_w_sum_one_range4302w(0);
	wire_man_prod_w_lg_w_vector1_range5228w5233w(0) <= wire_man_prod_w_vector1_range5228w(0) AND wire_man_prod_w_car_one_adj_range5227w(0);
	wire_man_prod_w_lg_w_vector1_range5228w5234w(0) <= wire_man_prod_w_vector1_range5228w(0) AND wire_man_prod_w_sum_one_range4312w(0);
	wire_man_prod_w_lg_w_vector1_range5239w5244w(0) <= wire_man_prod_w_vector1_range5239w(0) AND wire_man_prod_w_car_one_adj_range5238w(0);
	wire_man_prod_w_lg_w_vector1_range5239w5245w(0) <= wire_man_prod_w_vector1_range5239w(0) AND wire_man_prod_w_sum_one_range4322w(0);
	wire_man_prod_w_lg_w_vector1_range5250w5255w(0) <= wire_man_prod_w_vector1_range5250w(0) AND wire_man_prod_w_car_one_adj_range5249w(0);
	wire_man_prod_w_lg_w_vector1_range5250w5256w(0) <= wire_man_prod_w_vector1_range5250w(0) AND wire_man_prod_w_sum_one_range4332w(0);
	wire_man_prod_w_lg_w_vector1_range5261w5266w(0) <= wire_man_prod_w_vector1_range5261w(0) AND wire_man_prod_w_car_one_adj_range5260w(0);
	wire_man_prod_w_lg_w_vector1_range5261w5267w(0) <= wire_man_prod_w_vector1_range5261w(0) AND wire_man_prod_w_sum_one_range4342w(0);
	wire_man_prod_w_lg_w_vector1_range5272w5277w(0) <= wire_man_prod_w_vector1_range5272w(0) AND wire_man_prod_w_car_one_adj_range5271w(0);
	wire_man_prod_w_lg_w_vector1_range5272w5278w(0) <= wire_man_prod_w_vector1_range5272w(0) AND wire_man_prod_w_sum_one_range4352w(0);
	wire_man_prod_w_lg_w_vector1_range5283w5288w(0) <= wire_man_prod_w_vector1_range5283w(0) AND wire_man_prod_w_car_one_adj_range5282w(0);
	wire_man_prod_w_lg_w_vector1_range5283w5289w(0) <= wire_man_prod_w_vector1_range5283w(0) AND wire_man_prod_w_sum_one_range4362w(0);
	wire_man_prod_w_lg_w_vector1_range5294w5299w(0) <= wire_man_prod_w_vector1_range5294w(0) AND wire_man_prod_w_car_one_adj_range5293w(0);
	wire_man_prod_w_lg_w_vector1_range5294w5300w(0) <= wire_man_prod_w_vector1_range5294w(0) AND wire_man_prod_w_sum_one_range4372w(0);
	wire_man_prod_w_lg_w_vector1_range5305w5310w(0) <= wire_man_prod_w_vector1_range5305w(0) AND wire_man_prod_w_car_one_adj_range5304w(0);
	wire_man_prod_w_lg_w_vector1_range5305w5311w(0) <= wire_man_prod_w_vector1_range5305w(0) AND wire_man_prod_w_sum_one_range4382w(0);
	wire_man_prod_w_lg_w_vector1_range5107w5112w(0) <= wire_man_prod_w_vector1_range5107w(0) AND wire_man_prod_w_car_one_adj_range5106w(0);
	wire_man_prod_w_lg_w_vector1_range5107w5113w(0) <= wire_man_prod_w_vector1_range5107w(0) AND wire_man_prod_w_sum_one_range4202w(0);
	wire_man_prod_w_lg_w_vector1_range5316w5321w(0) <= wire_man_prod_w_vector1_range5316w(0) AND wire_man_prod_w_car_one_adj_range5315w(0);
	wire_man_prod_w_lg_w_vector1_range5316w5322w(0) <= wire_man_prod_w_vector1_range5316w(0) AND wire_man_prod_w_sum_one_range4392w(0);
	wire_man_prod_w_lg_w_vector1_range5327w5332w(0) <= wire_man_prod_w_vector1_range5327w(0) AND wire_man_prod_w_car_one_adj_range5326w(0);
	wire_man_prod_w_lg_w_vector1_range5327w5333w(0) <= wire_man_prod_w_vector1_range5327w(0) AND wire_man_prod_w_sum_one_range4402w(0);
	wire_man_prod_w_lg_w_vector1_range5338w5343w(0) <= wire_man_prod_w_vector1_range5338w(0) AND wire_man_prod_w_car_one_adj_range5337w(0);
	wire_man_prod_w_lg_w_vector1_range5338w5344w(0) <= wire_man_prod_w_vector1_range5338w(0) AND wire_man_prod_w_sum_one_range4412w(0);
	wire_man_prod_w_lg_w_vector1_range5349w5354w(0) <= wire_man_prod_w_vector1_range5349w(0) AND wire_man_prod_w_car_one_adj_range5348w(0);
	wire_man_prod_w_lg_w_vector1_range5349w5355w(0) <= wire_man_prod_w_vector1_range5349w(0) AND wire_man_prod_w_sum_one_range4422w(0);
	wire_man_prod_w_lg_w_vector1_range5360w5365w(0) <= wire_man_prod_w_vector1_range5360w(0) AND wire_man_prod_w_car_one_adj_range5359w(0);
	wire_man_prod_w_lg_w_vector1_range5360w5366w(0) <= wire_man_prod_w_vector1_range5360w(0) AND wire_man_prod_w_sum_one_range4432w(0);
	wire_man_prod_w_lg_w_vector1_range5371w5376w(0) <= wire_man_prod_w_vector1_range5371w(0) AND wire_man_prod_w_car_one_adj_range5370w(0);
	wire_man_prod_w_lg_w_vector1_range5371w5377w(0) <= wire_man_prod_w_vector1_range5371w(0) AND wire_man_prod_w_sum_one_range4442w(0);
	wire_man_prod_w_lg_w_vector1_range5382w5387w(0) <= wire_man_prod_w_vector1_range5382w(0) AND wire_man_prod_w_car_one_adj_range5381w(0);
	wire_man_prod_w_lg_w_vector1_range5382w5388w(0) <= wire_man_prod_w_vector1_range5382w(0) AND wire_man_prod_w_sum_one_range4452w(0);
	wire_man_prod_w_lg_w_vector1_range5393w5398w(0) <= wire_man_prod_w_vector1_range5393w(0) AND wire_man_prod_w_car_one_adj_range5392w(0);
	wire_man_prod_w_lg_w_vector1_range5393w5399w(0) <= wire_man_prod_w_vector1_range5393w(0) AND wire_man_prod_w_sum_one_range4462w(0);
	wire_man_prod_w_lg_w_vector1_range5404w5409w(0) <= wire_man_prod_w_vector1_range5404w(0) AND wire_man_prod_w_car_one_adj_range5403w(0);
	wire_man_prod_w_lg_w_vector1_range5404w5410w(0) <= wire_man_prod_w_vector1_range5404w(0) AND wire_man_prod_w_sum_one_range4472w(0);
	wire_man_prod_w_lg_w_vector1_range5415w5420w(0) <= wire_man_prod_w_vector1_range5415w(0) AND wire_man_prod_w_car_one_adj_range5414w(0);
	wire_man_prod_w_lg_w_vector1_range5415w5421w(0) <= wire_man_prod_w_vector1_range5415w(0) AND wire_man_prod_w_sum_one_range4482w(0);
	wire_man_prod_w_lg_w_vector1_range5118w5123w(0) <= wire_man_prod_w_vector1_range5118w(0) AND wire_man_prod_w_car_one_adj_range5117w(0);
	wire_man_prod_w_lg_w_vector1_range5118w5124w(0) <= wire_man_prod_w_vector1_range5118w(0) AND wire_man_prod_w_sum_one_range4212w(0);
	wire_man_prod_w_lg_w_vector1_range5426w5431w(0) <= wire_man_prod_w_vector1_range5426w(0) AND wire_man_prod_w_car_one_adj_range5425w(0);
	wire_man_prod_w_lg_w_vector1_range5426w5432w(0) <= wire_man_prod_w_vector1_range5426w(0) AND wire_man_prod_w_sum_one_range4492w(0);
	wire_man_prod_w_lg_w_vector1_range5437w5442w(0) <= wire_man_prod_w_vector1_range5437w(0) AND wire_man_prod_w_car_one_adj_range5436w(0);
	wire_man_prod_w_lg_w_vector1_range5437w5443w(0) <= wire_man_prod_w_vector1_range5437w(0) AND wire_man_prod_w_sum_one_range4502w(0);
	wire_man_prod_w_lg_w_vector1_range5448w5453w(0) <= wire_man_prod_w_vector1_range5448w(0) AND wire_man_prod_w_car_one_adj_range5447w(0);
	wire_man_prod_w_lg_w_vector1_range5448w5454w(0) <= wire_man_prod_w_vector1_range5448w(0) AND wire_man_prod_w_sum_one_range4512w(0);
	wire_man_prod_w_lg_w_vector1_range5459w5464w(0) <= wire_man_prod_w_vector1_range5459w(0) AND wire_man_prod_w_car_one_adj_range5458w(0);
	wire_man_prod_w_lg_w_vector1_range5459w5465w(0) <= wire_man_prod_w_vector1_range5459w(0) AND wire_man_prod_w_sum_one_range4522w(0);
	wire_man_prod_w_lg_w_vector1_range5470w5475w(0) <= wire_man_prod_w_vector1_range5470w(0) AND wire_man_prod_w_car_one_adj_range5469w(0);
	wire_man_prod_w_lg_w_vector1_range5470w5476w(0) <= wire_man_prod_w_vector1_range5470w(0) AND wire_man_prod_w_sum_one_range4532w(0);
	wire_man_prod_w_lg_w_vector1_range5481w5486w(0) <= wire_man_prod_w_vector1_range5481w(0) AND wire_man_prod_w_car_one_adj_range5480w(0);
	wire_man_prod_w_lg_w_vector1_range5481w5487w(0) <= wire_man_prod_w_vector1_range5481w(0) AND wire_man_prod_w_sum_one_range4542w(0);
	wire_man_prod_w_lg_w_vector1_range5492w5497w(0) <= wire_man_prod_w_vector1_range5492w(0) AND wire_man_prod_w_car_one_adj_range5491w(0);
	wire_man_prod_w_lg_w_vector1_range5492w5498w(0) <= wire_man_prod_w_vector1_range5492w(0) AND wire_man_prod_w_sum_one_range4552w(0);
	wire_man_prod_w_lg_w_vector1_range5503w5508w(0) <= wire_man_prod_w_vector1_range5503w(0) AND wire_man_prod_w_car_one_adj_range5502w(0);
	wire_man_prod_w_lg_w_vector1_range5503w5509w(0) <= wire_man_prod_w_vector1_range5503w(0) AND wire_man_prod_w_sum_one_range4562w(0);
	wire_man_prod_w_lg_w_vector1_range5514w5519w(0) <= wire_man_prod_w_vector1_range5514w(0) AND wire_man_prod_w_car_one_adj_range5513w(0);
	wire_man_prod_w_lg_w_vector1_range5514w5520w(0) <= wire_man_prod_w_vector1_range5514w(0) AND wire_man_prod_w_sum_one_range4572w(0);
	wire_man_prod_w_lg_w_vector1_range5525w5530w(0) <= wire_man_prod_w_vector1_range5525w(0) AND wire_man_prod_w_car_one_adj_range5524w(0);
	wire_man_prod_w_lg_w_vector1_range5525w5531w(0) <= wire_man_prod_w_vector1_range5525w(0) AND wire_man_prod_w_sum_one_range4582w(0);
	wire_man_prod_w_lg_w_vector1_range5129w5134w(0) <= wire_man_prod_w_vector1_range5129w(0) AND wire_man_prod_w_car_one_adj_range5128w(0);
	wire_man_prod_w_lg_w_vector1_range5129w5135w(0) <= wire_man_prod_w_vector1_range5129w(0) AND wire_man_prod_w_sum_one_range4222w(0);
	wire_man_prod_w_lg_w_vector1_range5536w5541w(0) <= wire_man_prod_w_vector1_range5536w(0) AND wire_man_prod_w_car_one_adj_range5535w(0);
	wire_man_prod_w_lg_w_vector1_range5536w5542w(0) <= wire_man_prod_w_vector1_range5536w(0) AND wire_man_prod_w_sum_one_range4592w(0);
	wire_man_prod_w_lg_w_vector1_range5547w5552w(0) <= wire_man_prod_w_vector1_range5547w(0) AND wire_man_prod_w_car_one_adj_range5546w(0);
	wire_man_prod_w_lg_w_vector1_range5547w5553w(0) <= wire_man_prod_w_vector1_range5547w(0) AND wire_man_prod_w_sum_one_range4602w(0);
	wire_man_prod_w_lg_w_vector1_range5558w5563w(0) <= wire_man_prod_w_vector1_range5558w(0) AND wire_man_prod_w_car_one_adj_range5557w(0);
	wire_man_prod_w_lg_w_vector1_range5558w5564w(0) <= wire_man_prod_w_vector1_range5558w(0) AND wire_man_prod_w_sum_one_range4612w(0);
	wire_man_prod_w_lg_w_vector1_range5569w5574w(0) <= wire_man_prod_w_vector1_range5569w(0) AND wire_man_prod_w_car_one_adj_range5568w(0);
	wire_man_prod_w_lg_w_vector1_range5569w5575w(0) <= wire_man_prod_w_vector1_range5569w(0) AND wire_man_prod_w_sum_one_range4622w(0);
	wire_man_prod_w_lg_w_vector1_range5580w5585w(0) <= wire_man_prod_w_vector1_range5580w(0) AND wire_man_prod_w_car_one_adj_range5579w(0);
	wire_man_prod_w_lg_w_vector1_range5580w5586w(0) <= wire_man_prod_w_vector1_range5580w(0) AND wire_man_prod_w_sum_one_range4632w(0);
	wire_man_prod_w_lg_w_vector1_range5591w5596w(0) <= wire_man_prod_w_vector1_range5591w(0) AND wire_man_prod_w_car_one_adj_range5590w(0);
	wire_man_prod_w_lg_w_vector1_range5591w5597w(0) <= wire_man_prod_w_vector1_range5591w(0) AND wire_man_prod_w_sum_one_range4642w(0);
	wire_man_prod_w_lg_w_vector1_range5602w5607w(0) <= wire_man_prod_w_vector1_range5602w(0) AND wire_man_prod_w_car_one_adj_range5601w(0);
	wire_man_prod_w_lg_w_vector1_range5602w5608w(0) <= wire_man_prod_w_vector1_range5602w(0) AND wire_man_prod_w_sum_one_range4652w(0);
	wire_man_prod_w_lg_w_vector1_range5613w5618w(0) <= wire_man_prod_w_vector1_range5613w(0) AND wire_man_prod_w_car_one_adj_range5612w(0);
	wire_man_prod_w_lg_w_vector1_range5613w5619w(0) <= wire_man_prod_w_vector1_range5613w(0) AND wire_man_prod_w_sum_one_range4662w(0);
	wire_man_prod_w_lg_w_vector1_range5624w5629w(0) <= wire_man_prod_w_vector1_range5624w(0) AND wire_man_prod_w_car_one_adj_range5623w(0);
	wire_man_prod_w_lg_w_vector1_range5624w5630w(0) <= wire_man_prod_w_vector1_range5624w(0) AND wire_man_prod_w_sum_one_range4672w(0);
	wire_man_prod_w_lg_w_vector1_range5635w5640w(0) <= wire_man_prod_w_vector1_range5635w(0) AND wire_man_prod_w_car_one_adj_range5634w(0);
	wire_man_prod_w_lg_w_vector1_range5635w5641w(0) <= wire_man_prod_w_vector1_range5635w(0) AND wire_man_prod_w_sum_one_range4682w(0);
	wire_man_prod_w_lg_w_vector1_range5140w5145w(0) <= wire_man_prod_w_vector1_range5140w(0) AND wire_man_prod_w_car_one_adj_range5139w(0);
	wire_man_prod_w_lg_w_vector1_range5140w5146w(0) <= wire_man_prod_w_vector1_range5140w(0) AND wire_man_prod_w_sum_one_range4232w(0);
	wire_man_prod_w_lg_w_vector1_range5646w5651w(0) <= wire_man_prod_w_vector1_range5646w(0) AND wire_man_prod_w_car_one_adj_range5645w(0);
	wire_man_prod_w_lg_w_vector1_range5646w5652w(0) <= wire_man_prod_w_vector1_range5646w(0) AND wire_man_prod_w_sum_one_range4692w(0);
	wire_man_prod_w_lg_w_vector1_range5657w5662w(0) <= wire_man_prod_w_vector1_range5657w(0) AND wire_man_prod_w_car_one_adj_range5656w(0);
	wire_man_prod_w_lg_w_vector1_range5657w5663w(0) <= wire_man_prod_w_vector1_range5657w(0) AND wire_man_prod_w_sum_one_range4702w(0);
	wire_man_prod_w_lg_w_vector1_range5668w5673w(0) <= wire_man_prod_w_vector1_range5668w(0) AND wire_man_prod_w_car_one_adj_range5667w(0);
	wire_man_prod_w_lg_w_vector1_range5668w5674w(0) <= wire_man_prod_w_vector1_range5668w(0) AND wire_man_prod_w_sum_one_range4712w(0);
	wire_man_prod_w_lg_w_vector1_range5679w5684w(0) <= wire_man_prod_w_vector1_range5679w(0) AND wire_man_prod_w_car_one_adj_range5678w(0);
	wire_man_prod_w_lg_w_vector1_range5679w5685w(0) <= wire_man_prod_w_vector1_range5679w(0) AND wire_man_prod_w_sum_one_range4722w(0);
	wire_man_prod_w_lg_w_vector1_range5690w5695w(0) <= wire_man_prod_w_vector1_range5690w(0) AND wire_man_prod_w_car_one_adj_range5689w(0);
	wire_man_prod_w_lg_w_vector1_range5690w5696w(0) <= wire_man_prod_w_vector1_range5690w(0) AND wire_man_prod_w_sum_one_range4732w(0);
	wire_man_prod_w_lg_w_vector1_range5701w5706w(0) <= wire_man_prod_w_vector1_range5701w(0) AND wire_man_prod_w_car_one_adj_range5700w(0);
	wire_man_prod_w_lg_w_vector1_range5701w5707w(0) <= wire_man_prod_w_vector1_range5701w(0) AND wire_man_prod_w_sum_one_range4742w(0);
	wire_man_prod_w_lg_w_vector1_range5712w5717w(0) <= wire_man_prod_w_vector1_range5712w(0) AND wire_man_prod_w_car_one_adj_range5711w(0);
	wire_man_prod_w_lg_w_vector1_range5712w5718w(0) <= wire_man_prod_w_vector1_range5712w(0) AND wire_man_prod_w_sum_one_range4752w(0);
	wire_man_prod_w_lg_w_vector1_range5723w5728w(0) <= wire_man_prod_w_vector1_range5723w(0) AND wire_man_prod_w_car_one_adj_range5722w(0);
	wire_man_prod_w_lg_w_vector1_range5723w5729w(0) <= wire_man_prod_w_vector1_range5723w(0) AND wire_man_prod_w_sum_one_range4762w(0);
	wire_man_prod_w_lg_w_vector1_range5734w5739w(0) <= wire_man_prod_w_vector1_range5734w(0) AND wire_man_prod_w_car_one_adj_range5733w(0);
	wire_man_prod_w_lg_w_vector1_range5734w5740w(0) <= wire_man_prod_w_vector1_range5734w(0) AND wire_man_prod_w_sum_one_range4772w(0);
	wire_man_prod_w_lg_w_vector1_range5745w5750w(0) <= wire_man_prod_w_vector1_range5745w(0) AND wire_man_prod_w_car_one_adj_range5744w(0);
	wire_man_prod_w_lg_w_vector1_range5745w5751w(0) <= wire_man_prod_w_vector1_range5745w(0) AND wire_man_prod_w_sum_one_range4782w(0);
	wire_man_prod_w_lg_w_vector1_range5151w5156w(0) <= wire_man_prod_w_vector1_range5151w(0) AND wire_man_prod_w_car_one_adj_range5150w(0);
	wire_man_prod_w_lg_w_vector1_range5151w5157w(0) <= wire_man_prod_w_vector1_range5151w(0) AND wire_man_prod_w_sum_one_range4242w(0);
	wire_man_prod_w_lg_w_vector1_range5756w5761w(0) <= wire_man_prod_w_vector1_range5756w(0) AND wire_man_prod_w_car_one_adj_range5755w(0);
	wire_man_prod_w_lg_w_vector1_range5756w5762w(0) <= wire_man_prod_w_vector1_range5756w(0) AND wire_man_prod_w_sum_one_range4792w(0);
	wire_man_prod_w_lg_w_vector1_range5767w5772w(0) <= wire_man_prod_w_vector1_range5767w(0) AND wire_man_prod_w_car_one_adj_range5766w(0);
	wire_man_prod_w_lg_w_vector1_range5767w5773w(0) <= wire_man_prod_w_vector1_range5767w(0) AND wire_man_prod_w_sum_one_range4802w(0);
	wire_man_prod_w_lg_w_vector1_range5778w5783w(0) <= wire_man_prod_w_vector1_range5778w(0) AND wire_man_prod_w_car_one_adj_range5777w(0);
	wire_man_prod_w_lg_w_vector1_range5778w5784w(0) <= wire_man_prod_w_vector1_range5778w(0) AND wire_man_prod_w_sum_one_range4812w(0);
	wire_man_prod_w_lg_w_vector1_range5789w5794w(0) <= wire_man_prod_w_vector1_range5789w(0) AND wire_man_prod_w_car_one_adj_range5788w(0);
	wire_man_prod_w_lg_w_vector1_range5789w5795w(0) <= wire_man_prod_w_vector1_range5789w(0) AND wire_man_prod_w_sum_one_range4822w(0);
	wire_man_prod_w_lg_w_vector1_range5800w5805w(0) <= wire_man_prod_w_vector1_range5800w(0) AND wire_man_prod_w_car_one_adj_range5799w(0);
	wire_man_prod_w_lg_w_vector1_range5800w5806w(0) <= wire_man_prod_w_vector1_range5800w(0) AND wire_man_prod_w_sum_one_range4832w(0);
	wire_man_prod_w_lg_w_vector1_range5811w5816w(0) <= wire_man_prod_w_vector1_range5811w(0) AND wire_man_prod_w_car_one_adj_range5810w(0);
	wire_man_prod_w_lg_w_vector1_range5811w5817w(0) <= wire_man_prod_w_vector1_range5811w(0) AND wire_man_prod_w_sum_one_range4842w(0);
	wire_man_prod_w_lg_w_vector1_range5822w5827w(0) <= wire_man_prod_w_vector1_range5822w(0) AND wire_man_prod_w_car_one_adj_range5821w(0);
	wire_man_prod_w_lg_w_vector1_range5822w5828w(0) <= wire_man_prod_w_vector1_range5822w(0) AND wire_man_prod_w_sum_one_range4852w(0);
	wire_man_prod_w_lg_w_vector1_range5833w5838w(0) <= wire_man_prod_w_vector1_range5833w(0) AND wire_man_prod_w_car_one_adj_range5832w(0);
	wire_man_prod_w_lg_w_vector1_range5833w5839w(0) <= wire_man_prod_w_vector1_range5833w(0) AND wire_man_prod_w_sum_one_range4862w(0);
	wire_man_prod_w_lg_w_vector1_range5844w5849w(0) <= wire_man_prod_w_vector1_range5844w(0) AND wire_man_prod_w_car_one_adj_range5843w(0);
	wire_man_prod_w_lg_w_vector1_range5844w5850w(0) <= wire_man_prod_w_vector1_range5844w(0) AND wire_man_prod_w_sum_one_range4872w(0);
	wire_man_prod_w_lg_w_vector1_range5855w5860w(0) <= wire_man_prod_w_vector1_range5855w(0) AND wire_man_prod_w_car_one_adj_range5854w(0);
	wire_man_prod_w_lg_w_vector1_range5855w5861w(0) <= wire_man_prod_w_vector1_range5855w(0) AND wire_man_prod_w_sum_one_range4882w(0);
	wire_man_prod_w_lg_w_vector1_range5162w5167w(0) <= wire_man_prod_w_vector1_range5162w(0) AND wire_man_prod_w_car_one_adj_range5161w(0);
	wire_man_prod_w_lg_w_vector1_range5162w5168w(0) <= wire_man_prod_w_vector1_range5162w(0) AND wire_man_prod_w_sum_one_range4252w(0);
	wire_man_prod_w_lg_w_vector1_range5866w5871w(0) <= wire_man_prod_w_vector1_range5866w(0) AND wire_man_prod_w_car_one_adj_range5865w(0);
	wire_man_prod_w_lg_w_vector1_range5866w5872w(0) <= wire_man_prod_w_vector1_range5866w(0) AND wire_man_prod_w_sum_one_range4892w(0);
	wire_man_prod_w_lg_w_vector1_range5877w5882w(0) <= wire_man_prod_w_vector1_range5877w(0) AND wire_man_prod_w_car_one_adj_range5876w(0);
	wire_man_prod_w_lg_w_vector1_range5877w5883w(0) <= wire_man_prod_w_vector1_range5877w(0) AND wire_man_prod_w_sum_one_range4902w(0);
	wire_man_prod_w_lg_w_vector1_range5888w5893w(0) <= wire_man_prod_w_vector1_range5888w(0) AND wire_man_prod_w_car_one_adj_range5887w(0);
	wire_man_prod_w_lg_w_vector1_range5888w5894w(0) <= wire_man_prod_w_vector1_range5888w(0) AND wire_man_prod_w_sum_one_range4912w(0);
	wire_man_prod_w_lg_w_vector1_range5899w5904w(0) <= wire_man_prod_w_vector1_range5899w(0) AND wire_man_prod_w_car_one_adj_range5898w(0);
	wire_man_prod_w_lg_w_vector1_range5899w5905w(0) <= wire_man_prod_w_vector1_range5899w(0) AND wire_man_prod_w_sum_one_range4922w(0);
	wire_man_prod_w_lg_w_vector1_range5910w5915w(0) <= wire_man_prod_w_vector1_range5910w(0) AND wire_man_prod_w_car_one_adj_range5909w(0);
	wire_man_prod_w_lg_w_vector1_range5910w5916w(0) <= wire_man_prod_w_vector1_range5910w(0) AND wire_man_prod_w_sum_one_range4932w(0);
	wire_man_prod_w_lg_w_vector1_range5921w5926w(0) <= wire_man_prod_w_vector1_range5921w(0) AND wire_man_prod_w_car_one_adj_range5920w(0);
	wire_man_prod_w_lg_w_vector1_range5921w5927w(0) <= wire_man_prod_w_vector1_range5921w(0) AND wire_man_prod_w_sum_one_range4942w(0);
	wire_man_prod_w_lg_w_vector1_range5932w5937w(0) <= wire_man_prod_w_vector1_range5932w(0) AND wire_man_prod_w_car_one_adj_range5931w(0);
	wire_man_prod_w_lg_w_vector1_range5932w5938w(0) <= wire_man_prod_w_vector1_range5932w(0) AND wire_man_prod_w_sum_one_range4952w(0);
	wire_man_prod_w_lg_w_vector1_range5943w5948w(0) <= wire_man_prod_w_vector1_range5943w(0) AND wire_man_prod_w_car_one_adj_range5942w(0);
	wire_man_prod_w_lg_w_vector1_range5943w5949w(0) <= wire_man_prod_w_vector1_range5943w(0) AND wire_man_prod_w_sum_one_range4962w(0);
	wire_man_prod_w_lg_w_vector1_range5954w5959w(0) <= wire_man_prod_w_vector1_range5954w(0) AND wire_man_prod_w_car_one_adj_range5953w(0);
	wire_man_prod_w_lg_w_vector1_range5954w5960w(0) <= wire_man_prod_w_vector1_range5954w(0) AND wire_man_prod_w_sum_one_range4972w(0);
	wire_man_prod_w_lg_w_vector1_range5965w5970w(0) <= wire_man_prod_w_vector1_range5965w(0) AND wire_man_prod_w_car_one_adj_range5964w(0);
	wire_man_prod_w_lg_w_vector1_range5965w5971w(0) <= wire_man_prod_w_vector1_range5965w(0) AND wire_man_prod_w_sum_one_range4982w(0);
	wire_man_prod_w_lg_w_vector1_range5173w5178w(0) <= wire_man_prod_w_vector1_range5173w(0) AND wire_man_prod_w_car_one_adj_range5172w(0);
	wire_man_prod_w_lg_w_vector1_range5173w5179w(0) <= wire_man_prod_w_vector1_range5173w(0) AND wire_man_prod_w_sum_one_range4262w(0);
	wire_man_prod_w_lg_w_vector1_range5976w5981w(0) <= wire_man_prod_w_vector1_range5976w(0) AND wire_man_prod_w_car_one_adj_range5975w(0);
	wire_man_prod_w_lg_w_vector1_range5976w5982w(0) <= wire_man_prod_w_vector1_range5976w(0) AND wire_man_prod_w_sum_one_range4992w(0);
	wire_man_prod_w_lg_w_vector1_range5987w5992w(0) <= wire_man_prod_w_vector1_range5987w(0) AND wire_man_prod_w_car_one_adj_range5986w(0);
	wire_man_prod_w_lg_w_vector1_range5987w5993w(0) <= wire_man_prod_w_vector1_range5987w(0) AND wire_man_prod_w_sum_one_range5002w(0);
	wire_man_prod_w_lg_w_vector1_range5998w6003w(0) <= wire_man_prod_w_vector1_range5998w(0) AND wire_man_prod_w_car_one_adj_range5997w(0);
	wire_man_prod_w_lg_w_vector1_range5998w6004w(0) <= wire_man_prod_w_vector1_range5998w(0) AND wire_man_prod_w_sum_one_range5012w(0);
	wire_man_prod_w_lg_w_vector1_range6009w6014w(0) <= wire_man_prod_w_vector1_range6009w(0) AND wire_man_prod_w_car_one_adj_range6008w(0);
	wire_man_prod_w_lg_w_vector1_range6009w6015w(0) <= wire_man_prod_w_vector1_range6009w(0) AND wire_man_prod_w_sum_one_range5022w(0);
	wire_man_prod_w_lg_w_vector1_range6020w6025w(0) <= wire_man_prod_w_vector1_range6020w(0) AND wire_man_prod_w_car_one_adj_range6019w(0);
	wire_man_prod_w_lg_w_vector1_range6020w6026w(0) <= wire_man_prod_w_vector1_range6020w(0) AND wire_man_prod_w_sum_one_range5032w(0);
	wire_man_prod_w_lg_w_vector1_range6031w6036w(0) <= wire_man_prod_w_vector1_range6031w(0) AND wire_man_prod_w_car_one_adj_range6030w(0);
	wire_man_prod_w_lg_w_vector1_range6031w6037w(0) <= wire_man_prod_w_vector1_range6031w(0) AND wire_man_prod_w_sum_one_range5042w(0);
	wire_man_prod_w_lg_w_vector1_range6042w6047w(0) <= wire_man_prod_w_vector1_range6042w(0) AND wire_man_prod_w_car_one_adj_range6041w(0);
	wire_man_prod_w_lg_w_vector1_range6042w6048w(0) <= wire_man_prod_w_vector1_range6042w(0) AND wire_man_prod_w_sum_one_range5052w(0);
	wire_man_prod_w_lg_w_vector1_range6053w6058w(0) <= wire_man_prod_w_vector1_range6053w(0) AND wire_man_prod_w_car_one_adj_range6052w(0);
	wire_man_prod_w_lg_w_vector1_range6053w6059w(0) <= wire_man_prod_w_vector1_range6053w(0) AND wire_man_prod_w_sum_one_range5062w(0);
	wire_man_prod_w_lg_w_vector1_range6064w6069w(0) <= wire_man_prod_w_vector1_range6064w(0) AND wire_man_prod_w_car_one_adj_range6063w(0);
	wire_man_prod_w_lg_w_vector1_range6064w6070w(0) <= wire_man_prod_w_vector1_range6064w(0) AND wire_man_prod_w_sum_one_range5072w(0);
	wire_man_prod_w_lg_w_vector1_range6075w6080w(0) <= wire_man_prod_w_vector1_range6075w(0) AND wire_man_prod_w_car_one_adj_range6074w(0);
	wire_man_prod_w_lg_w_vector1_range6075w6081w(0) <= wire_man_prod_w_vector1_range6075w(0) AND wire_man_prod_w_sum_one_range5082w(0);
	wire_man_prod_w_lg_w_vector1_range5184w5189w(0) <= wire_man_prod_w_vector1_range5184w(0) AND wire_man_prod_w_car_one_adj_range5183w(0);
	wire_man_prod_w_lg_w_vector1_range5184w5190w(0) <= wire_man_prod_w_vector1_range5184w(0) AND wire_man_prod_w_sum_one_range4272w(0);
	wire_man_prod_w_lg_w_vector1_range5195w5200w(0) <= wire_man_prod_w_vector1_range5195w(0) AND wire_man_prod_w_car_one_adj_range5194w(0);
	wire_man_prod_w_lg_w_vector1_range5195w5201w(0) <= wire_man_prod_w_vector1_range5195w(0) AND wire_man_prod_w_sum_one_range4282w(0);
	wire_man_prod_w_lg_w_vector2_range4187w4193w(0) <= wire_man_prod_w_vector2_range4187w(0) AND wire_man_prod_w_neg_lsb_range4186w(0);
	wire_man_prod_w_lg_w_vector2_range4187w4194w(0) <= wire_man_prod_w_vector2_range4187w(0) AND wire_man_prod_w_neg_msb_range4183w(0);
	wire_man_prod_w_lg_w_vector2_range4289w4294w(0) <= wire_man_prod_w_vector2_range4289w(0) AND wire_man_prod_w_neg_lsb_range4126w(0);
	wire_man_prod_w_lg_w_vector2_range4289w4295w(0) <= wire_man_prod_w_vector2_range4289w(0) AND wire_man_prod_w_neg_msb_range4123w(0);
	wire_man_prod_w_lg_w_vector2_range4299w4304w(0) <= wire_man_prod_w_vector2_range4299w(0) AND wire_man_prod_w_neg_lsb_range4120w(0);
	wire_man_prod_w_lg_w_vector2_range4299w4305w(0) <= wire_man_prod_w_vector2_range4299w(0) AND wire_man_prod_w_neg_msb_range4117w(0);
	wire_man_prod_w_lg_w_vector2_range4309w4314w(0) <= wire_man_prod_w_vector2_range4309w(0) AND wire_man_prod_w_neg_lsb_range4114w(0);
	wire_man_prod_w_lg_w_vector2_range4309w4315w(0) <= wire_man_prod_w_vector2_range4309w(0) AND wire_man_prod_w_neg_msb_range4111w(0);
	wire_man_prod_w_lg_w_vector2_range4319w4324w(0) <= wire_man_prod_w_vector2_range4319w(0) AND wire_man_prod_w_neg_lsb_range4108w(0);
	wire_man_prod_w_lg_w_vector2_range4319w4325w(0) <= wire_man_prod_w_vector2_range4319w(0) AND wire_man_prod_w_neg_msb_range4105w(0);
	wire_man_prod_w_lg_w_vector2_range4329w4334w(0) <= wire_man_prod_w_vector2_range4329w(0) AND wire_man_prod_w_neg_lsb_range4102w(0);
	wire_man_prod_w_lg_w_vector2_range4329w4335w(0) <= wire_man_prod_w_vector2_range4329w(0) AND wire_man_prod_w_neg_msb_range4099w(0);
	wire_man_prod_w_lg_w_vector2_range4339w4344w(0) <= wire_man_prod_w_vector2_range4339w(0) AND wire_man_prod_w_neg_lsb_range4096w(0);
	wire_man_prod_w_lg_w_vector2_range4339w4345w(0) <= wire_man_prod_w_vector2_range4339w(0) AND wire_man_prod_w_neg_msb_range4093w(0);
	wire_man_prod_w_lg_w_vector2_range4349w4354w(0) <= wire_man_prod_w_vector2_range4349w(0) AND wire_man_prod_w_neg_lsb_range4090w(0);
	wire_man_prod_w_lg_w_vector2_range4349w4355w(0) <= wire_man_prod_w_vector2_range4349w(0) AND wire_man_prod_w_neg_msb_range4087w(0);
	wire_man_prod_w_lg_w_vector2_range4359w4364w(0) <= wire_man_prod_w_vector2_range4359w(0) AND wire_man_prod_w_neg_lsb_range4084w(0);
	wire_man_prod_w_lg_w_vector2_range4359w4365w(0) <= wire_man_prod_w_vector2_range4359w(0) AND wire_man_prod_w_neg_msb_range4081w(0);
	wire_man_prod_w_lg_w_vector2_range4369w4374w(0) <= wire_man_prod_w_vector2_range4369w(0) AND wire_man_prod_w_neg_lsb_range4078w(0);
	wire_man_prod_w_lg_w_vector2_range4369w4375w(0) <= wire_man_prod_w_vector2_range4369w(0) AND wire_man_prod_w_neg_msb_range4075w(0);
	wire_man_prod_w_lg_w_vector2_range4379w4384w(0) <= wire_man_prod_w_vector2_range4379w(0) AND wire_man_prod_w_neg_lsb_range4072w(0);
	wire_man_prod_w_lg_w_vector2_range4379w4385w(0) <= wire_man_prod_w_vector2_range4379w(0) AND wire_man_prod_w_neg_msb_range4069w(0);
	wire_man_prod_w_lg_w_vector2_range4199w4204w(0) <= wire_man_prod_w_vector2_range4199w(0) AND wire_man_prod_w_neg_lsb_range4180w(0);
	wire_man_prod_w_lg_w_vector2_range4199w4205w(0) <= wire_man_prod_w_vector2_range4199w(0) AND wire_man_prod_w_neg_msb_range4177w(0);
	wire_man_prod_w_lg_w_vector2_range4389w4394w(0) <= wire_man_prod_w_vector2_range4389w(0) AND wire_man_prod_w_neg_lsb_range4066w(0);
	wire_man_prod_w_lg_w_vector2_range4389w4395w(0) <= wire_man_prod_w_vector2_range4389w(0) AND wire_man_prod_w_neg_msb_range4063w(0);
	wire_man_prod_w_lg_w_vector2_range4399w4404w(0) <= wire_man_prod_w_vector2_range4399w(0) AND wire_man_prod_w_neg_lsb_range4060w(0);
	wire_man_prod_w_lg_w_vector2_range4399w4405w(0) <= wire_man_prod_w_vector2_range4399w(0) AND wire_man_prod_w_neg_msb_range4057w(0);
	wire_man_prod_w_lg_w_vector2_range4409w4414w(0) <= wire_man_prod_w_vector2_range4409w(0) AND wire_man_prod_w_neg_lsb_range4054w(0);
	wire_man_prod_w_lg_w_vector2_range4409w4415w(0) <= wire_man_prod_w_vector2_range4409w(0) AND wire_man_prod_w_neg_msb_range4051w(0);
	wire_man_prod_w_lg_w_vector2_range4419w4424w(0) <= wire_man_prod_w_vector2_range4419w(0) AND wire_man_prod_w_neg_lsb_range4048w(0);
	wire_man_prod_w_lg_w_vector2_range4419w4425w(0) <= wire_man_prod_w_vector2_range4419w(0) AND wire_man_prod_w_neg_msb_range4045w(0);
	wire_man_prod_w_lg_w_vector2_range4429w4434w(0) <= wire_man_prod_w_vector2_range4429w(0) AND wire_man_prod_w_neg_lsb_range4042w(0);
	wire_man_prod_w_lg_w_vector2_range4429w4435w(0) <= wire_man_prod_w_vector2_range4429w(0) AND wire_man_prod_w_neg_msb_range4039w(0);
	wire_man_prod_w_lg_w_vector2_range4439w4444w(0) <= wire_man_prod_w_vector2_range4439w(0) AND wire_man_prod_w_neg_lsb_range4036w(0);
	wire_man_prod_w_lg_w_vector2_range4439w4445w(0) <= wire_man_prod_w_vector2_range4439w(0) AND wire_man_prod_w_neg_msb_range4033w(0);
	wire_man_prod_w_lg_w_vector2_range4449w4454w(0) <= wire_man_prod_w_vector2_range4449w(0) AND wire_man_prod_w_neg_lsb_range4030w(0);
	wire_man_prod_w_lg_w_vector2_range4449w4455w(0) <= wire_man_prod_w_vector2_range4449w(0) AND wire_man_prod_w_neg_msb_range4027w(0);
	wire_man_prod_w_lg_w_vector2_range4459w4464w(0) <= wire_man_prod_w_vector2_range4459w(0) AND wire_man_prod_w_neg_lsb_range4024w(0);
	wire_man_prod_w_lg_w_vector2_range4459w4465w(0) <= wire_man_prod_w_vector2_range4459w(0) AND wire_man_prod_w_neg_msb_range4021w(0);
	wire_man_prod_w_lg_w_vector2_range4469w4474w(0) <= wire_man_prod_w_vector2_range4469w(0) AND wire_man_prod_w_neg_lsb_range4018w(0);
	wire_man_prod_w_lg_w_vector2_range4469w4475w(0) <= wire_man_prod_w_vector2_range4469w(0) AND wire_man_prod_w_neg_msb_range4015w(0);
	wire_man_prod_w_lg_w_vector2_range4479w4484w(0) <= wire_man_prod_w_vector2_range4479w(0) AND wire_man_prod_w_neg_lsb_range4012w(0);
	wire_man_prod_w_lg_w_vector2_range4479w4485w(0) <= wire_man_prod_w_vector2_range4479w(0) AND wire_man_prod_w_neg_msb_range4009w(0);
	wire_man_prod_w_lg_w_vector2_range4209w4214w(0) <= wire_man_prod_w_vector2_range4209w(0) AND wire_man_prod_w_neg_lsb_range4174w(0);
	wire_man_prod_w_lg_w_vector2_range4209w4215w(0) <= wire_man_prod_w_vector2_range4209w(0) AND wire_man_prod_w_neg_msb_range4171w(0);
	wire_man_prod_w_lg_w_vector2_range4489w4494w(0) <= wire_man_prod_w_vector2_range4489w(0) AND wire_man_prod_w_neg_lsb_range4006w(0);
	wire_man_prod_w_lg_w_vector2_range4489w4495w(0) <= wire_man_prod_w_vector2_range4489w(0) AND wire_man_prod_w_neg_msb_range4003w(0);
	wire_man_prod_w_lg_w_vector2_range4499w4504w(0) <= wire_man_prod_w_vector2_range4499w(0) AND wire_man_prod_w_neg_lsb_range4000w(0);
	wire_man_prod_w_lg_w_vector2_range4499w4505w(0) <= wire_man_prod_w_vector2_range4499w(0) AND wire_man_prod_w_neg_msb_range3997w(0);
	wire_man_prod_w_lg_w_vector2_range4509w4514w(0) <= wire_man_prod_w_vector2_range4509w(0) AND wire_man_prod_w_neg_lsb_range3994w(0);
	wire_man_prod_w_lg_w_vector2_range4509w4515w(0) <= wire_man_prod_w_vector2_range4509w(0) AND wire_man_prod_w_neg_msb_range3991w(0);
	wire_man_prod_w_lg_w_vector2_range4519w4524w(0) <= wire_man_prod_w_vector2_range4519w(0) AND wire_man_prod_w_neg_lsb_range3988w(0);
	wire_man_prod_w_lg_w_vector2_range4519w4525w(0) <= wire_man_prod_w_vector2_range4519w(0) AND wire_man_prod_w_neg_msb_range3985w(0);
	wire_man_prod_w_lg_w_vector2_range4529w4534w(0) <= wire_man_prod_w_vector2_range4529w(0) AND wire_man_prod_w_neg_lsb_range3982w(0);
	wire_man_prod_w_lg_w_vector2_range4529w4535w(0) <= wire_man_prod_w_vector2_range4529w(0) AND wire_man_prod_w_neg_msb_range3979w(0);
	wire_man_prod_w_lg_w_vector2_range4539w4544w(0) <= wire_man_prod_w_vector2_range4539w(0) AND wire_man_prod_w_neg_lsb_range3976w(0);
	wire_man_prod_w_lg_w_vector2_range4539w4545w(0) <= wire_man_prod_w_vector2_range4539w(0) AND wire_man_prod_w_neg_msb_range3973w(0);
	wire_man_prod_w_lg_w_vector2_range4549w4554w(0) <= wire_man_prod_w_vector2_range4549w(0) AND wire_man_prod_w_neg_lsb_range3970w(0);
	wire_man_prod_w_lg_w_vector2_range4549w4555w(0) <= wire_man_prod_w_vector2_range4549w(0) AND wire_man_prod_w_neg_msb_range3967w(0);
	wire_man_prod_w_lg_w_vector2_range4559w4564w(0) <= wire_man_prod_w_vector2_range4559w(0) AND wire_man_prod_w_neg_lsb_range3964w(0);
	wire_man_prod_w_lg_w_vector2_range4559w4565w(0) <= wire_man_prod_w_vector2_range4559w(0) AND wire_man_prod_w_neg_msb_range3961w(0);
	wire_man_prod_w_lg_w_vector2_range4569w4574w(0) <= wire_man_prod_w_vector2_range4569w(0) AND wire_man_prod_w_neg_lsb_range3958w(0);
	wire_man_prod_w_lg_w_vector2_range4569w4575w(0) <= wire_man_prod_w_vector2_range4569w(0) AND wire_man_prod_w_neg_msb_range3955w(0);
	wire_man_prod_w_lg_w_vector2_range4579w4584w(0) <= wire_man_prod_w_vector2_range4579w(0) AND wire_man_prod_w_neg_lsb_range3952w(0);
	wire_man_prod_w_lg_w_vector2_range4579w4585w(0) <= wire_man_prod_w_vector2_range4579w(0) AND wire_man_prod_w_neg_msb_range3949w(0);
	wire_man_prod_w_lg_w_vector2_range4219w4224w(0) <= wire_man_prod_w_vector2_range4219w(0) AND wire_man_prod_w_neg_lsb_range4168w(0);
	wire_man_prod_w_lg_w_vector2_range4219w4225w(0) <= wire_man_prod_w_vector2_range4219w(0) AND wire_man_prod_w_neg_msb_range4165w(0);
	wire_man_prod_w_lg_w_vector2_range4589w4594w(0) <= wire_man_prod_w_vector2_range4589w(0) AND wire_man_prod_w_neg_lsb_range3946w(0);
	wire_man_prod_w_lg_w_vector2_range4589w4595w(0) <= wire_man_prod_w_vector2_range4589w(0) AND wire_man_prod_w_neg_msb_range3943w(0);
	wire_man_prod_w_lg_w_vector2_range4599w4604w(0) <= wire_man_prod_w_vector2_range4599w(0) AND wire_man_prod_w_neg_lsb_range3940w(0);
	wire_man_prod_w_lg_w_vector2_range4599w4605w(0) <= wire_man_prod_w_vector2_range4599w(0) AND wire_man_prod_w_neg_msb_range3937w(0);
	wire_man_prod_w_lg_w_vector2_range4609w4614w(0) <= wire_man_prod_w_vector2_range4609w(0) AND wire_man_prod_w_neg_lsb_range3934w(0);
	wire_man_prod_w_lg_w_vector2_range4609w4615w(0) <= wire_man_prod_w_vector2_range4609w(0) AND wire_man_prod_w_neg_msb_range3931w(0);
	wire_man_prod_w_lg_w_vector2_range4619w4624w(0) <= wire_man_prod_w_vector2_range4619w(0) AND wire_man_prod_w_neg_lsb_range3928w(0);
	wire_man_prod_w_lg_w_vector2_range4619w4625w(0) <= wire_man_prod_w_vector2_range4619w(0) AND wire_man_prod_w_neg_msb_range3925w(0);
	wire_man_prod_w_lg_w_vector2_range4629w4634w(0) <= wire_man_prod_w_vector2_range4629w(0) AND wire_man_prod_w_neg_lsb_range3922w(0);
	wire_man_prod_w_lg_w_vector2_range4629w4635w(0) <= wire_man_prod_w_vector2_range4629w(0) AND wire_man_prod_w_neg_msb_range3919w(0);
	wire_man_prod_w_lg_w_vector2_range4639w4644w(0) <= wire_man_prod_w_vector2_range4639w(0) AND wire_man_prod_w_neg_lsb_range3916w(0);
	wire_man_prod_w_lg_w_vector2_range4639w4645w(0) <= wire_man_prod_w_vector2_range4639w(0) AND wire_man_prod_w_neg_msb_range3913w(0);
	wire_man_prod_w_lg_w_vector2_range4649w4654w(0) <= wire_man_prod_w_vector2_range4649w(0) AND wire_man_prod_w_neg_lsb_range3910w(0);
	wire_man_prod_w_lg_w_vector2_range4649w4655w(0) <= wire_man_prod_w_vector2_range4649w(0) AND wire_man_prod_w_neg_msb_range3907w(0);
	wire_man_prod_w_lg_w_vector2_range4659w4664w(0) <= wire_man_prod_w_vector2_range4659w(0) AND wire_man_prod_w_neg_lsb_range3904w(0);
	wire_man_prod_w_lg_w_vector2_range4659w4665w(0) <= wire_man_prod_w_vector2_range4659w(0) AND wire_man_prod_w_neg_msb_range3901w(0);
	wire_man_prod_w_lg_w_vector2_range4669w4674w(0) <= wire_man_prod_w_vector2_range4669w(0) AND wire_man_prod_w_neg_lsb_range3898w(0);
	wire_man_prod_w_lg_w_vector2_range4669w4675w(0) <= wire_man_prod_w_vector2_range4669w(0) AND wire_man_prod_w_neg_msb_range3895w(0);
	wire_man_prod_w_lg_w_vector2_range4679w4684w(0) <= wire_man_prod_w_vector2_range4679w(0) AND wire_man_prod_w_neg_lsb_range3892w(0);
	wire_man_prod_w_lg_w_vector2_range4679w4685w(0) <= wire_man_prod_w_vector2_range4679w(0) AND wire_man_prod_w_neg_msb_range3889w(0);
	wire_man_prod_w_lg_w_vector2_range4229w4234w(0) <= wire_man_prod_w_vector2_range4229w(0) AND wire_man_prod_w_neg_lsb_range4162w(0);
	wire_man_prod_w_lg_w_vector2_range4229w4235w(0) <= wire_man_prod_w_vector2_range4229w(0) AND wire_man_prod_w_neg_msb_range4159w(0);
	wire_man_prod_w_lg_w_vector2_range4689w4694w(0) <= wire_man_prod_w_vector2_range4689w(0) AND wire_man_prod_w_neg_lsb_range3886w(0);
	wire_man_prod_w_lg_w_vector2_range4689w4695w(0) <= wire_man_prod_w_vector2_range4689w(0) AND wire_man_prod_w_neg_msb_range3883w(0);
	wire_man_prod_w_lg_w_vector2_range4699w4704w(0) <= wire_man_prod_w_vector2_range4699w(0) AND wire_man_prod_w_neg_lsb_range3880w(0);
	wire_man_prod_w_lg_w_vector2_range4699w4705w(0) <= wire_man_prod_w_vector2_range4699w(0) AND wire_man_prod_w_neg_msb_range3877w(0);
	wire_man_prod_w_lg_w_vector2_range4709w4714w(0) <= wire_man_prod_w_vector2_range4709w(0) AND wire_man_prod_w_neg_lsb_range3874w(0);
	wire_man_prod_w_lg_w_vector2_range4709w4715w(0) <= wire_man_prod_w_vector2_range4709w(0) AND wire_man_prod_w_neg_msb_range3871w(0);
	wire_man_prod_w_lg_w_vector2_range4719w4724w(0) <= wire_man_prod_w_vector2_range4719w(0) AND wire_man_prod_w_neg_lsb_range3868w(0);
	wire_man_prod_w_lg_w_vector2_range4719w4725w(0) <= wire_man_prod_w_vector2_range4719w(0) AND wire_man_prod_w_neg_msb_range3865w(0);
	wire_man_prod_w_lg_w_vector2_range4729w4734w(0) <= wire_man_prod_w_vector2_range4729w(0) AND wire_man_prod_w_neg_lsb_range3862w(0);
	wire_man_prod_w_lg_w_vector2_range4729w4735w(0) <= wire_man_prod_w_vector2_range4729w(0) AND wire_man_prod_w_neg_msb_range3859w(0);
	wire_man_prod_w_lg_w_vector2_range4739w4744w(0) <= wire_man_prod_w_vector2_range4739w(0) AND wire_man_prod_w_neg_lsb_range3856w(0);
	wire_man_prod_w_lg_w_vector2_range4739w4745w(0) <= wire_man_prod_w_vector2_range4739w(0) AND wire_man_prod_w_neg_msb_range3853w(0);
	wire_man_prod_w_lg_w_vector2_range4749w4754w(0) <= wire_man_prod_w_vector2_range4749w(0) AND wire_man_prod_w_neg_lsb_range3850w(0);
	wire_man_prod_w_lg_w_vector2_range4749w4755w(0) <= wire_man_prod_w_vector2_range4749w(0) AND wire_man_prod_w_neg_msb_range3847w(0);
	wire_man_prod_w_lg_w_vector2_range4759w4764w(0) <= wire_man_prod_w_vector2_range4759w(0) AND wire_man_prod_w_neg_lsb_range3844w(0);
	wire_man_prod_w_lg_w_vector2_range4759w4765w(0) <= wire_man_prod_w_vector2_range4759w(0) AND wire_man_prod_w_neg_msb_range3841w(0);
	wire_man_prod_w_lg_w_vector2_range4769w4774w(0) <= wire_man_prod_w_vector2_range4769w(0) AND wire_man_prod_w_neg_lsb_range3838w(0);
	wire_man_prod_w_lg_w_vector2_range4769w4775w(0) <= wire_man_prod_w_vector2_range4769w(0) AND wire_man_prod_w_neg_msb_range3835w(0);
	wire_man_prod_w_lg_w_vector2_range4779w4784w(0) <= wire_man_prod_w_vector2_range4779w(0) AND wire_man_prod_w_neg_lsb_range3832w(0);
	wire_man_prod_w_lg_w_vector2_range4779w4785w(0) <= wire_man_prod_w_vector2_range4779w(0) AND wire_man_prod_w_neg_msb_range3829w(0);
	wire_man_prod_w_lg_w_vector2_range4239w4244w(0) <= wire_man_prod_w_vector2_range4239w(0) AND wire_man_prod_w_neg_lsb_range4156w(0);
	wire_man_prod_w_lg_w_vector2_range4239w4245w(0) <= wire_man_prod_w_vector2_range4239w(0) AND wire_man_prod_w_neg_msb_range4153w(0);
	wire_man_prod_w_lg_w_vector2_range4789w4794w(0) <= wire_man_prod_w_vector2_range4789w(0) AND wire_man_prod_w_neg_lsb_range3825w(0);
	wire_man_prod_w_lg_w_vector2_range4789w4795w(0) <= wire_man_prod_w_vector2_range4789w(0) AND wire_man_prod_w_neg_msb_range3823w(0);
	wire_man_prod_w_lg_w_vector2_range4799w4804w(0) <= wire_man_prod_w_vector2_range4799w(0) AND wire_man_prod_w_neg_lsb_range3821w(0);
	wire_man_prod_w_lg_w_vector2_range4799w4805w(0) <= wire_man_prod_w_vector2_range4799w(0) AND wire_man_prod_w_neg_msb_range3819w(0);
	wire_man_prod_w_lg_w_vector2_range4809w4814w(0) <= wire_man_prod_w_vector2_range4809w(0) AND wire_man_prod_w_neg_lsb_range3817w(0);
	wire_man_prod_w_lg_w_vector2_range4809w4815w(0) <= wire_man_prod_w_vector2_range4809w(0) AND wire_man_prod_w_neg_msb_range3815w(0);
	wire_man_prod_w_lg_w_vector2_range4819w4824w(0) <= wire_man_prod_w_vector2_range4819w(0) AND wire_man_prod_w_neg_lsb_range3813w(0);
	wire_man_prod_w_lg_w_vector2_range4819w4825w(0) <= wire_man_prod_w_vector2_range4819w(0) AND wire_man_prod_w_neg_msb_range3811w(0);
	wire_man_prod_w_lg_w_vector2_range4829w4834w(0) <= wire_man_prod_w_vector2_range4829w(0) AND wire_man_prod_w_neg_lsb_range3809w(0);
	wire_man_prod_w_lg_w_vector2_range4829w4835w(0) <= wire_man_prod_w_vector2_range4829w(0) AND wire_man_prod_w_neg_msb_range3807w(0);
	wire_man_prod_w_lg_w_vector2_range4839w4844w(0) <= wire_man_prod_w_vector2_range4839w(0) AND wire_man_prod_w_neg_lsb_range3805w(0);
	wire_man_prod_w_lg_w_vector2_range4839w4845w(0) <= wire_man_prod_w_vector2_range4839w(0) AND wire_man_prod_w_neg_msb_range3803w(0);
	wire_man_prod_w_lg_w_vector2_range4849w4854w(0) <= wire_man_prod_w_vector2_range4849w(0) AND wire_man_prod_w_neg_lsb_range3801w(0);
	wire_man_prod_w_lg_w_vector2_range4849w4855w(0) <= wire_man_prod_w_vector2_range4849w(0) AND wire_man_prod_w_neg_msb_range3799w(0);
	wire_man_prod_w_lg_w_vector2_range4859w4864w(0) <= wire_man_prod_w_vector2_range4859w(0) AND wire_man_prod_w_neg_lsb_range3797w(0);
	wire_man_prod_w_lg_w_vector2_range4859w4865w(0) <= wire_man_prod_w_vector2_range4859w(0) AND wire_man_prod_w_neg_msb_range3795w(0);
	wire_man_prod_w_lg_w_vector2_range4869w4874w(0) <= wire_man_prod_w_vector2_range4869w(0) AND wire_man_prod_w_neg_lsb_range3793w(0);
	wire_man_prod_w_lg_w_vector2_range4869w4875w(0) <= wire_man_prod_w_vector2_range4869w(0) AND wire_man_prod_w_neg_msb_range3791w(0);
	wire_man_prod_w_lg_w_vector2_range4879w4884w(0) <= wire_man_prod_w_vector2_range4879w(0) AND wire_man_prod_w_neg_lsb_range3789w(0);
	wire_man_prod_w_lg_w_vector2_range4879w4885w(0) <= wire_man_prod_w_vector2_range4879w(0) AND wire_man_prod_w_neg_msb_range3787w(0);
	wire_man_prod_w_lg_w_vector2_range4249w4254w(0) <= wire_man_prod_w_vector2_range4249w(0) AND wire_man_prod_w_neg_lsb_range4150w(0);
	wire_man_prod_w_lg_w_vector2_range4249w4255w(0) <= wire_man_prod_w_vector2_range4249w(0) AND wire_man_prod_w_neg_msb_range4147w(0);
	wire_man_prod_w_lg_w_vector2_range4889w4894w(0) <= wire_man_prod_w_vector2_range4889w(0) AND wire_man_prod_w_neg_lsb_range3785w(0);
	wire_man_prod_w_lg_w_vector2_range4889w4895w(0) <= wire_man_prod_w_vector2_range4889w(0) AND wire_man_prod_w_neg_msb_range3783w(0);
	wire_man_prod_w_lg_w_vector2_range4899w4904w(0) <= wire_man_prod_w_vector2_range4899w(0) AND wire_man_prod_w_neg_lsb_range3781w(0);
	wire_man_prod_w_lg_w_vector2_range4899w4905w(0) <= wire_man_prod_w_vector2_range4899w(0) AND wire_man_prod_w_neg_msb_range3779w(0);
	wire_man_prod_w_lg_w_vector2_range4909w4914w(0) <= wire_man_prod_w_vector2_range4909w(0) AND wire_man_prod_w_neg_lsb_range3777w(0);
	wire_man_prod_w_lg_w_vector2_range4909w4915w(0) <= wire_man_prod_w_vector2_range4909w(0) AND wire_man_prod_w_neg_msb_range3775w(0);
	wire_man_prod_w_lg_w_vector2_range4919w4924w(0) <= wire_man_prod_w_vector2_range4919w(0) AND wire_man_prod_w_neg_lsb_range3773w(0);
	wire_man_prod_w_lg_w_vector2_range4919w4925w(0) <= wire_man_prod_w_vector2_range4919w(0) AND wire_man_prod_w_neg_msb_range3771w(0);
	wire_man_prod_w_lg_w_vector2_range4929w4934w(0) <= wire_man_prod_w_vector2_range4929w(0) AND wire_man_prod_w_neg_lsb_range3769w(0);
	wire_man_prod_w_lg_w_vector2_range4929w4935w(0) <= wire_man_prod_w_vector2_range4929w(0) AND wire_man_prod_w_neg_msb_range3767w(0);
	wire_man_prod_w_lg_w_vector2_range4939w4944w(0) <= wire_man_prod_w_vector2_range4939w(0) AND wire_man_prod_w_neg_lsb_range3765w(0);
	wire_man_prod_w_lg_w_vector2_range4939w4945w(0) <= wire_man_prod_w_vector2_range4939w(0) AND wire_man_prod_w_neg_msb_range3763w(0);
	wire_man_prod_w_lg_w_vector2_range4949w4954w(0) <= wire_man_prod_w_vector2_range4949w(0) AND wire_man_prod_w_neg_lsb_range3761w(0);
	wire_man_prod_w_lg_w_vector2_range4949w4955w(0) <= wire_man_prod_w_vector2_range4949w(0) AND wire_man_prod_w_neg_msb_range3759w(0);
	wire_man_prod_w_lg_w_vector2_range4959w4964w(0) <= wire_man_prod_w_vector2_range4959w(0) AND wire_man_prod_w_neg_lsb_range3757w(0);
	wire_man_prod_w_lg_w_vector2_range4959w4965w(0) <= wire_man_prod_w_vector2_range4959w(0) AND wire_man_prod_w_neg_msb_range3755w(0);
	wire_man_prod_w_lg_w_vector2_range4969w4974w(0) <= wire_man_prod_w_vector2_range4969w(0) AND wire_man_prod_w_neg_lsb_range3753w(0);
	wire_man_prod_w_lg_w_vector2_range4969w4975w(0) <= wire_man_prod_w_vector2_range4969w(0) AND wire_man_prod_w_neg_msb_range3751w(0);
	wire_man_prod_w_lg_w_vector2_range4979w4984w(0) <= wire_man_prod_w_vector2_range4979w(0) AND wire_man_prod_w_neg_lsb_range3749w(0);
	wire_man_prod_w_lg_w_vector2_range4979w4985w(0) <= wire_man_prod_w_vector2_range4979w(0) AND wire_man_prod_w_neg_msb_range3747w(0);
	wire_man_prod_w_lg_w_vector2_range4259w4264w(0) <= wire_man_prod_w_vector2_range4259w(0) AND wire_man_prod_w_neg_lsb_range4144w(0);
	wire_man_prod_w_lg_w_vector2_range4259w4265w(0) <= wire_man_prod_w_vector2_range4259w(0) AND wire_man_prod_w_neg_msb_range4141w(0);
	wire_man_prod_w_lg_w_vector2_range4989w4994w(0) <= wire_man_prod_w_vector2_range4989w(0) AND wire_man_prod_w_neg_lsb_range3745w(0);
	wire_man_prod_w_lg_w_vector2_range4989w4995w(0) <= wire_man_prod_w_vector2_range4989w(0) AND wire_man_prod_w_neg_msb_range3743w(0);
	wire_man_prod_w_lg_w_vector2_range4999w5004w(0) <= wire_man_prod_w_vector2_range4999w(0) AND wire_man_prod_w_neg_lsb_range3741w(0);
	wire_man_prod_w_lg_w_vector2_range4999w5005w(0) <= wire_man_prod_w_vector2_range4999w(0) AND wire_man_prod_w_neg_msb_range3739w(0);
	wire_man_prod_w_lg_w_vector2_range5009w5014w(0) <= wire_man_prod_w_vector2_range5009w(0) AND wire_man_prod_w_neg_lsb_range3737w(0);
	wire_man_prod_w_lg_w_vector2_range5009w5015w(0) <= wire_man_prod_w_vector2_range5009w(0) AND wire_man_prod_w_neg_msb_range3735w(0);
	wire_man_prod_w_lg_w_vector2_range5019w5024w(0) <= wire_man_prod_w_vector2_range5019w(0) AND wire_man_prod_w_neg_lsb_range3733w(0);
	wire_man_prod_w_lg_w_vector2_range5019w5025w(0) <= wire_man_prod_w_vector2_range5019w(0) AND wire_man_prod_w_neg_msb_range3731w(0);
	wire_man_prod_w_lg_w_vector2_range5029w5034w(0) <= wire_man_prod_w_vector2_range5029w(0) AND wire_man_prod_w_neg_lsb_range3729w(0);
	wire_man_prod_w_lg_w_vector2_range5029w5035w(0) <= wire_man_prod_w_vector2_range5029w(0) AND wire_man_prod_w_neg_msb_range3727w(0);
	wire_man_prod_w_lg_w_vector2_range5039w5044w(0) <= wire_man_prod_w_vector2_range5039w(0) AND wire_man_prod_w_neg_lsb_range3725w(0);
	wire_man_prod_w_lg_w_vector2_range5039w5045w(0) <= wire_man_prod_w_vector2_range5039w(0) AND wire_man_prod_w_neg_msb_range3723w(0);
	wire_man_prod_w_lg_w_vector2_range5049w5054w(0) <= wire_man_prod_w_vector2_range5049w(0) AND wire_man_prod_w_neg_lsb_range3721w(0);
	wire_man_prod_w_lg_w_vector2_range5049w5055w(0) <= wire_man_prod_w_vector2_range5049w(0) AND wire_man_prod_w_neg_msb_range3719w(0);
	wire_man_prod_w_lg_w_vector2_range5059w5064w(0) <= wire_man_prod_w_vector2_range5059w(0) AND wire_man_prod_w_neg_lsb_range3717w(0);
	wire_man_prod_w_lg_w_vector2_range5059w5065w(0) <= wire_man_prod_w_vector2_range5059w(0) AND wire_man_prod_w_neg_msb_range3715w(0);
	wire_man_prod_w_lg_w_vector2_range5069w5074w(0) <= wire_man_prod_w_vector2_range5069w(0) AND wire_man_prod_w_neg_lsb_range3713w(0);
	wire_man_prod_w_lg_w_vector2_range5069w5075w(0) <= wire_man_prod_w_vector2_range5069w(0) AND wire_man_prod_w_neg_msb_range3711w(0);
	wire_man_prod_w_lg_w_vector2_range5079w5084w(0) <= wire_man_prod_w_vector2_range5079w(0) AND wire_man_prod_w_neg_lsb_range3708w(0);
	wire_man_prod_w_lg_w_vector2_range5079w5085w(0) <= wire_man_prod_w_vector2_range5079w(0) AND wire_man_prod_w_neg_msb_range3705w(0);
	wire_man_prod_w_lg_w_vector2_range4269w4274w(0) <= wire_man_prod_w_vector2_range4269w(0) AND wire_man_prod_w_neg_lsb_range4138w(0);
	wire_man_prod_w_lg_w_vector2_range4269w4275w(0) <= wire_man_prod_w_vector2_range4269w(0) AND wire_man_prod_w_neg_msb_range4135w(0);
	wire_man_prod_w_lg_w_vector2_range4279w4284w(0) <= wire_man_prod_w_vector2_range4279w(0) AND wire_man_prod_w_neg_lsb_range4132w(0);
	wire_man_prod_w_lg_w_vector2_range4279w4285w(0) <= wire_man_prod_w_vector2_range4279w(0) AND wire_man_prod_w_neg_msb_range4129w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4184w4185w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4184w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4124w4125w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4124w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4118w4119w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4118w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4112w4113w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4112w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4106w4107w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4106w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4100w4101w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4100w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4094w4095w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4094w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4088w4089w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4088w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4082w4083w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4082w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4076w4077w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4076w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4070w4071w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4070w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4178w4179w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4178w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4064w4065w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4064w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4058w4059w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4058w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4052w4053w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4052w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4046w4047w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4046w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4040w4041w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4040w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4034w4035w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4034w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4028w4029w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4028w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4022w4023w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4022w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4016w4017w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4016w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4010w4011w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4010w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4172w4173w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4172w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4004w4005w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4004w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3998w3999w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3998w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3992w3993w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3992w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3986w3987w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3986w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3980w3981w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3980w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3974w3975w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3974w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3968w3969w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3968w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3962w3963w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3962w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3956w3957w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3956w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3950w3951w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3950w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4166w4167w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4166w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3944w3945w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3944w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3938w3939w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3938w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3932w3933w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3932w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3926w3927w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3926w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3920w3921w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3920w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3914w3915w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3914w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3908w3909w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3908w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3902w3903w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3902w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3896w3897w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3896w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3890w3891w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3890w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4160w4161w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4160w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3884w3885w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3884w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3878w3879w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3878w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3872w3873w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3872w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3866w3867w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3866w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3860w3861w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3860w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3854w3855w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3854w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3848w3849w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3848w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3842w3843w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3842w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3836w3837w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3836w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range3830w3831w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range3830w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4154w4155w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4154w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4148w4149w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4148w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4142w4143w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4142w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4136w4137w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4136w(0);
	wire_man_prod_w_lg_w_lsb_prod_wo_range4130w4131w(0) <= NOT wire_man_prod_w_lsb_prod_wo_range4130w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4181w4182w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4181w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4121w4122w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4121w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4115w4116w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4115w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4109w4110w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4109w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4103w4104w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4103w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4097w4098w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4097w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4091w4092w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4091w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4085w4086w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4085w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4079w4080w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4079w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4073w4074w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4073w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4067w4068w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4067w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4175w4176w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4175w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4061w4062w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4061w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4055w4056w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4055w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4049w4050w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4049w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4043w4044w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4043w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4037w4038w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4037w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4031w4032w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4031w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4025w4026w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4025w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4019w4020w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4019w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4013w4014w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4013w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4007w4008w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4007w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4169w4170w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4169w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4001w4002w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4001w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3995w3996w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3995w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3989w3990w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3989w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3983w3984w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3983w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3977w3978w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3977w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3971w3972w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3971w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3965w3966w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3965w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3959w3960w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3959w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3953w3954w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3953w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3947w3948w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3947w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4163w4164w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4163w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3941w3942w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3941w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3935w3936w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3935w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3929w3930w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3929w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3923w3924w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3923w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3917w3918w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3917w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3911w3912w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3911w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3905w3906w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3905w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3899w3900w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3899w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3893w3894w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3893w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3887w3888w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3887w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4157w4158w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4157w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3881w3882w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3881w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3875w3876w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3875w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3869w3870w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3869w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3863w3864w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3863w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3857w3858w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3857w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3851w3852w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3851w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3845w3846w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3845w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3839w3840w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3839w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3833w3834w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3833w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range3827w3828w(0) <= NOT wire_man_prod_w_msb_prod_wo_range3827w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4151w4152w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4151w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4145w4146w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4145w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4139w4140w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4139w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4133w4134w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4133w(0);
	wire_man_prod_w_lg_w_msb_prod_wo_range4127w4128w(0) <= NOT wire_man_prod_w_msb_prod_wo_range4127w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5094w5101w5102w(0) <= wire_man_prod_w_lg_w_vector1_range5094w5101w(0) OR wire_man_prod_w_lg_w_vector1_range5094w5100w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5206w5212w5213w(0) <= wire_man_prod_w_lg_w_vector1_range5206w5212w(0) OR wire_man_prod_w_lg_w_vector1_range5206w5211w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5217w5223w5224w(0) <= wire_man_prod_w_lg_w_vector1_range5217w5223w(0) OR wire_man_prod_w_lg_w_vector1_range5217w5222w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5228w5234w5235w(0) <= wire_man_prod_w_lg_w_vector1_range5228w5234w(0) OR wire_man_prod_w_lg_w_vector1_range5228w5233w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5239w5245w5246w(0) <= wire_man_prod_w_lg_w_vector1_range5239w5245w(0) OR wire_man_prod_w_lg_w_vector1_range5239w5244w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5250w5256w5257w(0) <= wire_man_prod_w_lg_w_vector1_range5250w5256w(0) OR wire_man_prod_w_lg_w_vector1_range5250w5255w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5261w5267w5268w(0) <= wire_man_prod_w_lg_w_vector1_range5261w5267w(0) OR wire_man_prod_w_lg_w_vector1_range5261w5266w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5272w5278w5279w(0) <= wire_man_prod_w_lg_w_vector1_range5272w5278w(0) OR wire_man_prod_w_lg_w_vector1_range5272w5277w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5283w5289w5290w(0) <= wire_man_prod_w_lg_w_vector1_range5283w5289w(0) OR wire_man_prod_w_lg_w_vector1_range5283w5288w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5294w5300w5301w(0) <= wire_man_prod_w_lg_w_vector1_range5294w5300w(0) OR wire_man_prod_w_lg_w_vector1_range5294w5299w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5305w5311w5312w(0) <= wire_man_prod_w_lg_w_vector1_range5305w5311w(0) OR wire_man_prod_w_lg_w_vector1_range5305w5310w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5107w5113w5114w(0) <= wire_man_prod_w_lg_w_vector1_range5107w5113w(0) OR wire_man_prod_w_lg_w_vector1_range5107w5112w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5316w5322w5323w(0) <= wire_man_prod_w_lg_w_vector1_range5316w5322w(0) OR wire_man_prod_w_lg_w_vector1_range5316w5321w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5327w5333w5334w(0) <= wire_man_prod_w_lg_w_vector1_range5327w5333w(0) OR wire_man_prod_w_lg_w_vector1_range5327w5332w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5338w5344w5345w(0) <= wire_man_prod_w_lg_w_vector1_range5338w5344w(0) OR wire_man_prod_w_lg_w_vector1_range5338w5343w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5349w5355w5356w(0) <= wire_man_prod_w_lg_w_vector1_range5349w5355w(0) OR wire_man_prod_w_lg_w_vector1_range5349w5354w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5360w5366w5367w(0) <= wire_man_prod_w_lg_w_vector1_range5360w5366w(0) OR wire_man_prod_w_lg_w_vector1_range5360w5365w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5371w5377w5378w(0) <= wire_man_prod_w_lg_w_vector1_range5371w5377w(0) OR wire_man_prod_w_lg_w_vector1_range5371w5376w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5382w5388w5389w(0) <= wire_man_prod_w_lg_w_vector1_range5382w5388w(0) OR wire_man_prod_w_lg_w_vector1_range5382w5387w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5393w5399w5400w(0) <= wire_man_prod_w_lg_w_vector1_range5393w5399w(0) OR wire_man_prod_w_lg_w_vector1_range5393w5398w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5404w5410w5411w(0) <= wire_man_prod_w_lg_w_vector1_range5404w5410w(0) OR wire_man_prod_w_lg_w_vector1_range5404w5409w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5415w5421w5422w(0) <= wire_man_prod_w_lg_w_vector1_range5415w5421w(0) OR wire_man_prod_w_lg_w_vector1_range5415w5420w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5118w5124w5125w(0) <= wire_man_prod_w_lg_w_vector1_range5118w5124w(0) OR wire_man_prod_w_lg_w_vector1_range5118w5123w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5426w5432w5433w(0) <= wire_man_prod_w_lg_w_vector1_range5426w5432w(0) OR wire_man_prod_w_lg_w_vector1_range5426w5431w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5437w5443w5444w(0) <= wire_man_prod_w_lg_w_vector1_range5437w5443w(0) OR wire_man_prod_w_lg_w_vector1_range5437w5442w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5448w5454w5455w(0) <= wire_man_prod_w_lg_w_vector1_range5448w5454w(0) OR wire_man_prod_w_lg_w_vector1_range5448w5453w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5459w5465w5466w(0) <= wire_man_prod_w_lg_w_vector1_range5459w5465w(0) OR wire_man_prod_w_lg_w_vector1_range5459w5464w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5470w5476w5477w(0) <= wire_man_prod_w_lg_w_vector1_range5470w5476w(0) OR wire_man_prod_w_lg_w_vector1_range5470w5475w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5481w5487w5488w(0) <= wire_man_prod_w_lg_w_vector1_range5481w5487w(0) OR wire_man_prod_w_lg_w_vector1_range5481w5486w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5492w5498w5499w(0) <= wire_man_prod_w_lg_w_vector1_range5492w5498w(0) OR wire_man_prod_w_lg_w_vector1_range5492w5497w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5503w5509w5510w(0) <= wire_man_prod_w_lg_w_vector1_range5503w5509w(0) OR wire_man_prod_w_lg_w_vector1_range5503w5508w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5514w5520w5521w(0) <= wire_man_prod_w_lg_w_vector1_range5514w5520w(0) OR wire_man_prod_w_lg_w_vector1_range5514w5519w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5525w5531w5532w(0) <= wire_man_prod_w_lg_w_vector1_range5525w5531w(0) OR wire_man_prod_w_lg_w_vector1_range5525w5530w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5129w5135w5136w(0) <= wire_man_prod_w_lg_w_vector1_range5129w5135w(0) OR wire_man_prod_w_lg_w_vector1_range5129w5134w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5536w5542w5543w(0) <= wire_man_prod_w_lg_w_vector1_range5536w5542w(0) OR wire_man_prod_w_lg_w_vector1_range5536w5541w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5547w5553w5554w(0) <= wire_man_prod_w_lg_w_vector1_range5547w5553w(0) OR wire_man_prod_w_lg_w_vector1_range5547w5552w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5558w5564w5565w(0) <= wire_man_prod_w_lg_w_vector1_range5558w5564w(0) OR wire_man_prod_w_lg_w_vector1_range5558w5563w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5569w5575w5576w(0) <= wire_man_prod_w_lg_w_vector1_range5569w5575w(0) OR wire_man_prod_w_lg_w_vector1_range5569w5574w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5580w5586w5587w(0) <= wire_man_prod_w_lg_w_vector1_range5580w5586w(0) OR wire_man_prod_w_lg_w_vector1_range5580w5585w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5591w5597w5598w(0) <= wire_man_prod_w_lg_w_vector1_range5591w5597w(0) OR wire_man_prod_w_lg_w_vector1_range5591w5596w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5602w5608w5609w(0) <= wire_man_prod_w_lg_w_vector1_range5602w5608w(0) OR wire_man_prod_w_lg_w_vector1_range5602w5607w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5613w5619w5620w(0) <= wire_man_prod_w_lg_w_vector1_range5613w5619w(0) OR wire_man_prod_w_lg_w_vector1_range5613w5618w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5624w5630w5631w(0) <= wire_man_prod_w_lg_w_vector1_range5624w5630w(0) OR wire_man_prod_w_lg_w_vector1_range5624w5629w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5635w5641w5642w(0) <= wire_man_prod_w_lg_w_vector1_range5635w5641w(0) OR wire_man_prod_w_lg_w_vector1_range5635w5640w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5140w5146w5147w(0) <= wire_man_prod_w_lg_w_vector1_range5140w5146w(0) OR wire_man_prod_w_lg_w_vector1_range5140w5145w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5646w5652w5653w(0) <= wire_man_prod_w_lg_w_vector1_range5646w5652w(0) OR wire_man_prod_w_lg_w_vector1_range5646w5651w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5657w5663w5664w(0) <= wire_man_prod_w_lg_w_vector1_range5657w5663w(0) OR wire_man_prod_w_lg_w_vector1_range5657w5662w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5668w5674w5675w(0) <= wire_man_prod_w_lg_w_vector1_range5668w5674w(0) OR wire_man_prod_w_lg_w_vector1_range5668w5673w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5679w5685w5686w(0) <= wire_man_prod_w_lg_w_vector1_range5679w5685w(0) OR wire_man_prod_w_lg_w_vector1_range5679w5684w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5690w5696w5697w(0) <= wire_man_prod_w_lg_w_vector1_range5690w5696w(0) OR wire_man_prod_w_lg_w_vector1_range5690w5695w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5701w5707w5708w(0) <= wire_man_prod_w_lg_w_vector1_range5701w5707w(0) OR wire_man_prod_w_lg_w_vector1_range5701w5706w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5712w5718w5719w(0) <= wire_man_prod_w_lg_w_vector1_range5712w5718w(0) OR wire_man_prod_w_lg_w_vector1_range5712w5717w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5723w5729w5730w(0) <= wire_man_prod_w_lg_w_vector1_range5723w5729w(0) OR wire_man_prod_w_lg_w_vector1_range5723w5728w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5734w5740w5741w(0) <= wire_man_prod_w_lg_w_vector1_range5734w5740w(0) OR wire_man_prod_w_lg_w_vector1_range5734w5739w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5745w5751w5752w(0) <= wire_man_prod_w_lg_w_vector1_range5745w5751w(0) OR wire_man_prod_w_lg_w_vector1_range5745w5750w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5151w5157w5158w(0) <= wire_man_prod_w_lg_w_vector1_range5151w5157w(0) OR wire_man_prod_w_lg_w_vector1_range5151w5156w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5756w5762w5763w(0) <= wire_man_prod_w_lg_w_vector1_range5756w5762w(0) OR wire_man_prod_w_lg_w_vector1_range5756w5761w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5767w5773w5774w(0) <= wire_man_prod_w_lg_w_vector1_range5767w5773w(0) OR wire_man_prod_w_lg_w_vector1_range5767w5772w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5778w5784w5785w(0) <= wire_man_prod_w_lg_w_vector1_range5778w5784w(0) OR wire_man_prod_w_lg_w_vector1_range5778w5783w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5789w5795w5796w(0) <= wire_man_prod_w_lg_w_vector1_range5789w5795w(0) OR wire_man_prod_w_lg_w_vector1_range5789w5794w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5800w5806w5807w(0) <= wire_man_prod_w_lg_w_vector1_range5800w5806w(0) OR wire_man_prod_w_lg_w_vector1_range5800w5805w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5811w5817w5818w(0) <= wire_man_prod_w_lg_w_vector1_range5811w5817w(0) OR wire_man_prod_w_lg_w_vector1_range5811w5816w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5822w5828w5829w(0) <= wire_man_prod_w_lg_w_vector1_range5822w5828w(0) OR wire_man_prod_w_lg_w_vector1_range5822w5827w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5833w5839w5840w(0) <= wire_man_prod_w_lg_w_vector1_range5833w5839w(0) OR wire_man_prod_w_lg_w_vector1_range5833w5838w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5844w5850w5851w(0) <= wire_man_prod_w_lg_w_vector1_range5844w5850w(0) OR wire_man_prod_w_lg_w_vector1_range5844w5849w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5855w5861w5862w(0) <= wire_man_prod_w_lg_w_vector1_range5855w5861w(0) OR wire_man_prod_w_lg_w_vector1_range5855w5860w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5162w5168w5169w(0) <= wire_man_prod_w_lg_w_vector1_range5162w5168w(0) OR wire_man_prod_w_lg_w_vector1_range5162w5167w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5866w5872w5873w(0) <= wire_man_prod_w_lg_w_vector1_range5866w5872w(0) OR wire_man_prod_w_lg_w_vector1_range5866w5871w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5877w5883w5884w(0) <= wire_man_prod_w_lg_w_vector1_range5877w5883w(0) OR wire_man_prod_w_lg_w_vector1_range5877w5882w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5888w5894w5895w(0) <= wire_man_prod_w_lg_w_vector1_range5888w5894w(0) OR wire_man_prod_w_lg_w_vector1_range5888w5893w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5899w5905w5906w(0) <= wire_man_prod_w_lg_w_vector1_range5899w5905w(0) OR wire_man_prod_w_lg_w_vector1_range5899w5904w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5910w5916w5917w(0) <= wire_man_prod_w_lg_w_vector1_range5910w5916w(0) OR wire_man_prod_w_lg_w_vector1_range5910w5915w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5921w5927w5928w(0) <= wire_man_prod_w_lg_w_vector1_range5921w5927w(0) OR wire_man_prod_w_lg_w_vector1_range5921w5926w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5932w5938w5939w(0) <= wire_man_prod_w_lg_w_vector1_range5932w5938w(0) OR wire_man_prod_w_lg_w_vector1_range5932w5937w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5943w5949w5950w(0) <= wire_man_prod_w_lg_w_vector1_range5943w5949w(0) OR wire_man_prod_w_lg_w_vector1_range5943w5948w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5954w5960w5961w(0) <= wire_man_prod_w_lg_w_vector1_range5954w5960w(0) OR wire_man_prod_w_lg_w_vector1_range5954w5959w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5965w5971w5972w(0) <= wire_man_prod_w_lg_w_vector1_range5965w5971w(0) OR wire_man_prod_w_lg_w_vector1_range5965w5970w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5173w5179w5180w(0) <= wire_man_prod_w_lg_w_vector1_range5173w5179w(0) OR wire_man_prod_w_lg_w_vector1_range5173w5178w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5976w5982w5983w(0) <= wire_man_prod_w_lg_w_vector1_range5976w5982w(0) OR wire_man_prod_w_lg_w_vector1_range5976w5981w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5987w5993w5994w(0) <= wire_man_prod_w_lg_w_vector1_range5987w5993w(0) OR wire_man_prod_w_lg_w_vector1_range5987w5992w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5998w6004w6005w(0) <= wire_man_prod_w_lg_w_vector1_range5998w6004w(0) OR wire_man_prod_w_lg_w_vector1_range5998w6003w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6009w6015w6016w(0) <= wire_man_prod_w_lg_w_vector1_range6009w6015w(0) OR wire_man_prod_w_lg_w_vector1_range6009w6014w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6020w6026w6027w(0) <= wire_man_prod_w_lg_w_vector1_range6020w6026w(0) OR wire_man_prod_w_lg_w_vector1_range6020w6025w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6031w6037w6038w(0) <= wire_man_prod_w_lg_w_vector1_range6031w6037w(0) OR wire_man_prod_w_lg_w_vector1_range6031w6036w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6042w6048w6049w(0) <= wire_man_prod_w_lg_w_vector1_range6042w6048w(0) OR wire_man_prod_w_lg_w_vector1_range6042w6047w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6053w6059w6060w(0) <= wire_man_prod_w_lg_w_vector1_range6053w6059w(0) OR wire_man_prod_w_lg_w_vector1_range6053w6058w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6064w6070w6071w(0) <= wire_man_prod_w_lg_w_vector1_range6064w6070w(0) OR wire_man_prod_w_lg_w_vector1_range6064w6069w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6075w6081w6082w(0) <= wire_man_prod_w_lg_w_vector1_range6075w6081w(0) OR wire_man_prod_w_lg_w_vector1_range6075w6080w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5184w5190w5191w(0) <= wire_man_prod_w_lg_w_vector1_range5184w5190w(0) OR wire_man_prod_w_lg_w_vector1_range5184w5189w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5195w5201w5202w(0) <= wire_man_prod_w_lg_w_vector1_range5195w5201w(0) OR wire_man_prod_w_lg_w_vector1_range5195w5200w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4187w4194w4195w(0) <= wire_man_prod_w_lg_w_vector2_range4187w4194w(0) OR wire_man_prod_w_lg_w_vector2_range4187w4193w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4289w4295w4296w(0) <= wire_man_prod_w_lg_w_vector2_range4289w4295w(0) OR wire_man_prod_w_lg_w_vector2_range4289w4294w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4299w4305w4306w(0) <= wire_man_prod_w_lg_w_vector2_range4299w4305w(0) OR wire_man_prod_w_lg_w_vector2_range4299w4304w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4309w4315w4316w(0) <= wire_man_prod_w_lg_w_vector2_range4309w4315w(0) OR wire_man_prod_w_lg_w_vector2_range4309w4314w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4319w4325w4326w(0) <= wire_man_prod_w_lg_w_vector2_range4319w4325w(0) OR wire_man_prod_w_lg_w_vector2_range4319w4324w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4329w4335w4336w(0) <= wire_man_prod_w_lg_w_vector2_range4329w4335w(0) OR wire_man_prod_w_lg_w_vector2_range4329w4334w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4339w4345w4346w(0) <= wire_man_prod_w_lg_w_vector2_range4339w4345w(0) OR wire_man_prod_w_lg_w_vector2_range4339w4344w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4349w4355w4356w(0) <= wire_man_prod_w_lg_w_vector2_range4349w4355w(0) OR wire_man_prod_w_lg_w_vector2_range4349w4354w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4359w4365w4366w(0) <= wire_man_prod_w_lg_w_vector2_range4359w4365w(0) OR wire_man_prod_w_lg_w_vector2_range4359w4364w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4369w4375w4376w(0) <= wire_man_prod_w_lg_w_vector2_range4369w4375w(0) OR wire_man_prod_w_lg_w_vector2_range4369w4374w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4379w4385w4386w(0) <= wire_man_prod_w_lg_w_vector2_range4379w4385w(0) OR wire_man_prod_w_lg_w_vector2_range4379w4384w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4199w4205w4206w(0) <= wire_man_prod_w_lg_w_vector2_range4199w4205w(0) OR wire_man_prod_w_lg_w_vector2_range4199w4204w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4389w4395w4396w(0) <= wire_man_prod_w_lg_w_vector2_range4389w4395w(0) OR wire_man_prod_w_lg_w_vector2_range4389w4394w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4399w4405w4406w(0) <= wire_man_prod_w_lg_w_vector2_range4399w4405w(0) OR wire_man_prod_w_lg_w_vector2_range4399w4404w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4409w4415w4416w(0) <= wire_man_prod_w_lg_w_vector2_range4409w4415w(0) OR wire_man_prod_w_lg_w_vector2_range4409w4414w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4419w4425w4426w(0) <= wire_man_prod_w_lg_w_vector2_range4419w4425w(0) OR wire_man_prod_w_lg_w_vector2_range4419w4424w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4429w4435w4436w(0) <= wire_man_prod_w_lg_w_vector2_range4429w4435w(0) OR wire_man_prod_w_lg_w_vector2_range4429w4434w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4439w4445w4446w(0) <= wire_man_prod_w_lg_w_vector2_range4439w4445w(0) OR wire_man_prod_w_lg_w_vector2_range4439w4444w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4449w4455w4456w(0) <= wire_man_prod_w_lg_w_vector2_range4449w4455w(0) OR wire_man_prod_w_lg_w_vector2_range4449w4454w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4459w4465w4466w(0) <= wire_man_prod_w_lg_w_vector2_range4459w4465w(0) OR wire_man_prod_w_lg_w_vector2_range4459w4464w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4469w4475w4476w(0) <= wire_man_prod_w_lg_w_vector2_range4469w4475w(0) OR wire_man_prod_w_lg_w_vector2_range4469w4474w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4479w4485w4486w(0) <= wire_man_prod_w_lg_w_vector2_range4479w4485w(0) OR wire_man_prod_w_lg_w_vector2_range4479w4484w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4209w4215w4216w(0) <= wire_man_prod_w_lg_w_vector2_range4209w4215w(0) OR wire_man_prod_w_lg_w_vector2_range4209w4214w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4489w4495w4496w(0) <= wire_man_prod_w_lg_w_vector2_range4489w4495w(0) OR wire_man_prod_w_lg_w_vector2_range4489w4494w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4499w4505w4506w(0) <= wire_man_prod_w_lg_w_vector2_range4499w4505w(0) OR wire_man_prod_w_lg_w_vector2_range4499w4504w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4509w4515w4516w(0) <= wire_man_prod_w_lg_w_vector2_range4509w4515w(0) OR wire_man_prod_w_lg_w_vector2_range4509w4514w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4519w4525w4526w(0) <= wire_man_prod_w_lg_w_vector2_range4519w4525w(0) OR wire_man_prod_w_lg_w_vector2_range4519w4524w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4529w4535w4536w(0) <= wire_man_prod_w_lg_w_vector2_range4529w4535w(0) OR wire_man_prod_w_lg_w_vector2_range4529w4534w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4539w4545w4546w(0) <= wire_man_prod_w_lg_w_vector2_range4539w4545w(0) OR wire_man_prod_w_lg_w_vector2_range4539w4544w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4549w4555w4556w(0) <= wire_man_prod_w_lg_w_vector2_range4549w4555w(0) OR wire_man_prod_w_lg_w_vector2_range4549w4554w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4559w4565w4566w(0) <= wire_man_prod_w_lg_w_vector2_range4559w4565w(0) OR wire_man_prod_w_lg_w_vector2_range4559w4564w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4569w4575w4576w(0) <= wire_man_prod_w_lg_w_vector2_range4569w4575w(0) OR wire_man_prod_w_lg_w_vector2_range4569w4574w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4579w4585w4586w(0) <= wire_man_prod_w_lg_w_vector2_range4579w4585w(0) OR wire_man_prod_w_lg_w_vector2_range4579w4584w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4219w4225w4226w(0) <= wire_man_prod_w_lg_w_vector2_range4219w4225w(0) OR wire_man_prod_w_lg_w_vector2_range4219w4224w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4589w4595w4596w(0) <= wire_man_prod_w_lg_w_vector2_range4589w4595w(0) OR wire_man_prod_w_lg_w_vector2_range4589w4594w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4599w4605w4606w(0) <= wire_man_prod_w_lg_w_vector2_range4599w4605w(0) OR wire_man_prod_w_lg_w_vector2_range4599w4604w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4609w4615w4616w(0) <= wire_man_prod_w_lg_w_vector2_range4609w4615w(0) OR wire_man_prod_w_lg_w_vector2_range4609w4614w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4619w4625w4626w(0) <= wire_man_prod_w_lg_w_vector2_range4619w4625w(0) OR wire_man_prod_w_lg_w_vector2_range4619w4624w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4629w4635w4636w(0) <= wire_man_prod_w_lg_w_vector2_range4629w4635w(0) OR wire_man_prod_w_lg_w_vector2_range4629w4634w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4639w4645w4646w(0) <= wire_man_prod_w_lg_w_vector2_range4639w4645w(0) OR wire_man_prod_w_lg_w_vector2_range4639w4644w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4649w4655w4656w(0) <= wire_man_prod_w_lg_w_vector2_range4649w4655w(0) OR wire_man_prod_w_lg_w_vector2_range4649w4654w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4659w4665w4666w(0) <= wire_man_prod_w_lg_w_vector2_range4659w4665w(0) OR wire_man_prod_w_lg_w_vector2_range4659w4664w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4669w4675w4676w(0) <= wire_man_prod_w_lg_w_vector2_range4669w4675w(0) OR wire_man_prod_w_lg_w_vector2_range4669w4674w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4679w4685w4686w(0) <= wire_man_prod_w_lg_w_vector2_range4679w4685w(0) OR wire_man_prod_w_lg_w_vector2_range4679w4684w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4229w4235w4236w(0) <= wire_man_prod_w_lg_w_vector2_range4229w4235w(0) OR wire_man_prod_w_lg_w_vector2_range4229w4234w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4689w4695w4696w(0) <= wire_man_prod_w_lg_w_vector2_range4689w4695w(0) OR wire_man_prod_w_lg_w_vector2_range4689w4694w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4699w4705w4706w(0) <= wire_man_prod_w_lg_w_vector2_range4699w4705w(0) OR wire_man_prod_w_lg_w_vector2_range4699w4704w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4709w4715w4716w(0) <= wire_man_prod_w_lg_w_vector2_range4709w4715w(0) OR wire_man_prod_w_lg_w_vector2_range4709w4714w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4719w4725w4726w(0) <= wire_man_prod_w_lg_w_vector2_range4719w4725w(0) OR wire_man_prod_w_lg_w_vector2_range4719w4724w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4729w4735w4736w(0) <= wire_man_prod_w_lg_w_vector2_range4729w4735w(0) OR wire_man_prod_w_lg_w_vector2_range4729w4734w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4739w4745w4746w(0) <= wire_man_prod_w_lg_w_vector2_range4739w4745w(0) OR wire_man_prod_w_lg_w_vector2_range4739w4744w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4749w4755w4756w(0) <= wire_man_prod_w_lg_w_vector2_range4749w4755w(0) OR wire_man_prod_w_lg_w_vector2_range4749w4754w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4759w4765w4766w(0) <= wire_man_prod_w_lg_w_vector2_range4759w4765w(0) OR wire_man_prod_w_lg_w_vector2_range4759w4764w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4769w4775w4776w(0) <= wire_man_prod_w_lg_w_vector2_range4769w4775w(0) OR wire_man_prod_w_lg_w_vector2_range4769w4774w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4779w4785w4786w(0) <= wire_man_prod_w_lg_w_vector2_range4779w4785w(0) OR wire_man_prod_w_lg_w_vector2_range4779w4784w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4239w4245w4246w(0) <= wire_man_prod_w_lg_w_vector2_range4239w4245w(0) OR wire_man_prod_w_lg_w_vector2_range4239w4244w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4789w4795w4796w(0) <= wire_man_prod_w_lg_w_vector2_range4789w4795w(0) OR wire_man_prod_w_lg_w_vector2_range4789w4794w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4799w4805w4806w(0) <= wire_man_prod_w_lg_w_vector2_range4799w4805w(0) OR wire_man_prod_w_lg_w_vector2_range4799w4804w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4809w4815w4816w(0) <= wire_man_prod_w_lg_w_vector2_range4809w4815w(0) OR wire_man_prod_w_lg_w_vector2_range4809w4814w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4819w4825w4826w(0) <= wire_man_prod_w_lg_w_vector2_range4819w4825w(0) OR wire_man_prod_w_lg_w_vector2_range4819w4824w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4829w4835w4836w(0) <= wire_man_prod_w_lg_w_vector2_range4829w4835w(0) OR wire_man_prod_w_lg_w_vector2_range4829w4834w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4839w4845w4846w(0) <= wire_man_prod_w_lg_w_vector2_range4839w4845w(0) OR wire_man_prod_w_lg_w_vector2_range4839w4844w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4849w4855w4856w(0) <= wire_man_prod_w_lg_w_vector2_range4849w4855w(0) OR wire_man_prod_w_lg_w_vector2_range4849w4854w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4859w4865w4866w(0) <= wire_man_prod_w_lg_w_vector2_range4859w4865w(0) OR wire_man_prod_w_lg_w_vector2_range4859w4864w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4869w4875w4876w(0) <= wire_man_prod_w_lg_w_vector2_range4869w4875w(0) OR wire_man_prod_w_lg_w_vector2_range4869w4874w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4879w4885w4886w(0) <= wire_man_prod_w_lg_w_vector2_range4879w4885w(0) OR wire_man_prod_w_lg_w_vector2_range4879w4884w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4249w4255w4256w(0) <= wire_man_prod_w_lg_w_vector2_range4249w4255w(0) OR wire_man_prod_w_lg_w_vector2_range4249w4254w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4889w4895w4896w(0) <= wire_man_prod_w_lg_w_vector2_range4889w4895w(0) OR wire_man_prod_w_lg_w_vector2_range4889w4894w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4899w4905w4906w(0) <= wire_man_prod_w_lg_w_vector2_range4899w4905w(0) OR wire_man_prod_w_lg_w_vector2_range4899w4904w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4909w4915w4916w(0) <= wire_man_prod_w_lg_w_vector2_range4909w4915w(0) OR wire_man_prod_w_lg_w_vector2_range4909w4914w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4919w4925w4926w(0) <= wire_man_prod_w_lg_w_vector2_range4919w4925w(0) OR wire_man_prod_w_lg_w_vector2_range4919w4924w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4929w4935w4936w(0) <= wire_man_prod_w_lg_w_vector2_range4929w4935w(0) OR wire_man_prod_w_lg_w_vector2_range4929w4934w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4939w4945w4946w(0) <= wire_man_prod_w_lg_w_vector2_range4939w4945w(0) OR wire_man_prod_w_lg_w_vector2_range4939w4944w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4949w4955w4956w(0) <= wire_man_prod_w_lg_w_vector2_range4949w4955w(0) OR wire_man_prod_w_lg_w_vector2_range4949w4954w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4959w4965w4966w(0) <= wire_man_prod_w_lg_w_vector2_range4959w4965w(0) OR wire_man_prod_w_lg_w_vector2_range4959w4964w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4969w4975w4976w(0) <= wire_man_prod_w_lg_w_vector2_range4969w4975w(0) OR wire_man_prod_w_lg_w_vector2_range4969w4974w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4979w4985w4986w(0) <= wire_man_prod_w_lg_w_vector2_range4979w4985w(0) OR wire_man_prod_w_lg_w_vector2_range4979w4984w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4259w4265w4266w(0) <= wire_man_prod_w_lg_w_vector2_range4259w4265w(0) OR wire_man_prod_w_lg_w_vector2_range4259w4264w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4989w4995w4996w(0) <= wire_man_prod_w_lg_w_vector2_range4989w4995w(0) OR wire_man_prod_w_lg_w_vector2_range4989w4994w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4999w5005w5006w(0) <= wire_man_prod_w_lg_w_vector2_range4999w5005w(0) OR wire_man_prod_w_lg_w_vector2_range4999w5004w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5009w5015w5016w(0) <= wire_man_prod_w_lg_w_vector2_range5009w5015w(0) OR wire_man_prod_w_lg_w_vector2_range5009w5014w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5019w5025w5026w(0) <= wire_man_prod_w_lg_w_vector2_range5019w5025w(0) OR wire_man_prod_w_lg_w_vector2_range5019w5024w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5029w5035w5036w(0) <= wire_man_prod_w_lg_w_vector2_range5029w5035w(0) OR wire_man_prod_w_lg_w_vector2_range5029w5034w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5039w5045w5046w(0) <= wire_man_prod_w_lg_w_vector2_range5039w5045w(0) OR wire_man_prod_w_lg_w_vector2_range5039w5044w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5049w5055w5056w(0) <= wire_man_prod_w_lg_w_vector2_range5049w5055w(0) OR wire_man_prod_w_lg_w_vector2_range5049w5054w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5059w5065w5066w(0) <= wire_man_prod_w_lg_w_vector2_range5059w5065w(0) OR wire_man_prod_w_lg_w_vector2_range5059w5064w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5069w5075w5076w(0) <= wire_man_prod_w_lg_w_vector2_range5069w5075w(0) OR wire_man_prod_w_lg_w_vector2_range5069w5074w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5079w5085w5086w(0) <= wire_man_prod_w_lg_w_vector2_range5079w5085w(0) OR wire_man_prod_w_lg_w_vector2_range5079w5084w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4269w4275w4276w(0) <= wire_man_prod_w_lg_w_vector2_range4269w4275w(0) OR wire_man_prod_w_lg_w_vector2_range4269w4274w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4279w4285w4286w(0) <= wire_man_prod_w_lg_w_vector2_range4279w4285w(0) OR wire_man_prod_w_lg_w_vector2_range4279w4284w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5094w5101w5102w5103w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5094w5101w5102w(0) OR wire_man_prod_w_lg_w_sum_one_range4190w5099w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5206w5212w5213w5214w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5206w5212w5213w(0) OR wire_man_prod_w_lg_w_sum_one_range4292w5210w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5217w5223w5224w5225w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5217w5223w5224w(0) OR wire_man_prod_w_lg_w_sum_one_range4302w5221w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5228w5234w5235w5236w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5228w5234w5235w(0) OR wire_man_prod_w_lg_w_sum_one_range4312w5232w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5239w5245w5246w5247w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5239w5245w5246w(0) OR wire_man_prod_w_lg_w_sum_one_range4322w5243w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5250w5256w5257w5258w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5250w5256w5257w(0) OR wire_man_prod_w_lg_w_sum_one_range4332w5254w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5261w5267w5268w5269w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5261w5267w5268w(0) OR wire_man_prod_w_lg_w_sum_one_range4342w5265w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5272w5278w5279w5280w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5272w5278w5279w(0) OR wire_man_prod_w_lg_w_sum_one_range4352w5276w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5283w5289w5290w5291w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5283w5289w5290w(0) OR wire_man_prod_w_lg_w_sum_one_range4362w5287w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5294w5300w5301w5302w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5294w5300w5301w(0) OR wire_man_prod_w_lg_w_sum_one_range4372w5298w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5305w5311w5312w5313w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5305w5311w5312w(0) OR wire_man_prod_w_lg_w_sum_one_range4382w5309w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5107w5113w5114w5115w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5107w5113w5114w(0) OR wire_man_prod_w_lg_w_sum_one_range4202w5111w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5316w5322w5323w5324w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5316w5322w5323w(0) OR wire_man_prod_w_lg_w_sum_one_range4392w5320w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5327w5333w5334w5335w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5327w5333w5334w(0) OR wire_man_prod_w_lg_w_sum_one_range4402w5331w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5338w5344w5345w5346w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5338w5344w5345w(0) OR wire_man_prod_w_lg_w_sum_one_range4412w5342w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5349w5355w5356w5357w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5349w5355w5356w(0) OR wire_man_prod_w_lg_w_sum_one_range4422w5353w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5360w5366w5367w5368w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5360w5366w5367w(0) OR wire_man_prod_w_lg_w_sum_one_range4432w5364w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5371w5377w5378w5379w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5371w5377w5378w(0) OR wire_man_prod_w_lg_w_sum_one_range4442w5375w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5382w5388w5389w5390w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5382w5388w5389w(0) OR wire_man_prod_w_lg_w_sum_one_range4452w5386w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5393w5399w5400w5401w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5393w5399w5400w(0) OR wire_man_prod_w_lg_w_sum_one_range4462w5397w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5404w5410w5411w5412w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5404w5410w5411w(0) OR wire_man_prod_w_lg_w_sum_one_range4472w5408w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5415w5421w5422w5423w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5415w5421w5422w(0) OR wire_man_prod_w_lg_w_sum_one_range4482w5419w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5118w5124w5125w5126w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5118w5124w5125w(0) OR wire_man_prod_w_lg_w_sum_one_range4212w5122w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5426w5432w5433w5434w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5426w5432w5433w(0) OR wire_man_prod_w_lg_w_sum_one_range4492w5430w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5437w5443w5444w5445w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5437w5443w5444w(0) OR wire_man_prod_w_lg_w_sum_one_range4502w5441w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5448w5454w5455w5456w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5448w5454w5455w(0) OR wire_man_prod_w_lg_w_sum_one_range4512w5452w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5459w5465w5466w5467w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5459w5465w5466w(0) OR wire_man_prod_w_lg_w_sum_one_range4522w5463w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5470w5476w5477w5478w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5470w5476w5477w(0) OR wire_man_prod_w_lg_w_sum_one_range4532w5474w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5481w5487w5488w5489w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5481w5487w5488w(0) OR wire_man_prod_w_lg_w_sum_one_range4542w5485w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5492w5498w5499w5500w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5492w5498w5499w(0) OR wire_man_prod_w_lg_w_sum_one_range4552w5496w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5503w5509w5510w5511w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5503w5509w5510w(0) OR wire_man_prod_w_lg_w_sum_one_range4562w5507w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5514w5520w5521w5522w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5514w5520w5521w(0) OR wire_man_prod_w_lg_w_sum_one_range4572w5518w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5525w5531w5532w5533w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5525w5531w5532w(0) OR wire_man_prod_w_lg_w_sum_one_range4582w5529w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5129w5135w5136w5137w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5129w5135w5136w(0) OR wire_man_prod_w_lg_w_sum_one_range4222w5133w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5536w5542w5543w5544w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5536w5542w5543w(0) OR wire_man_prod_w_lg_w_sum_one_range4592w5540w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5547w5553w5554w5555w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5547w5553w5554w(0) OR wire_man_prod_w_lg_w_sum_one_range4602w5551w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5558w5564w5565w5566w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5558w5564w5565w(0) OR wire_man_prod_w_lg_w_sum_one_range4612w5562w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5569w5575w5576w5577w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5569w5575w5576w(0) OR wire_man_prod_w_lg_w_sum_one_range4622w5573w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5580w5586w5587w5588w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5580w5586w5587w(0) OR wire_man_prod_w_lg_w_sum_one_range4632w5584w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5591w5597w5598w5599w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5591w5597w5598w(0) OR wire_man_prod_w_lg_w_sum_one_range4642w5595w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5602w5608w5609w5610w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5602w5608w5609w(0) OR wire_man_prod_w_lg_w_sum_one_range4652w5606w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5613w5619w5620w5621w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5613w5619w5620w(0) OR wire_man_prod_w_lg_w_sum_one_range4662w5617w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5624w5630w5631w5632w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5624w5630w5631w(0) OR wire_man_prod_w_lg_w_sum_one_range4672w5628w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5635w5641w5642w5643w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5635w5641w5642w(0) OR wire_man_prod_w_lg_w_sum_one_range4682w5639w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5140w5146w5147w5148w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5140w5146w5147w(0) OR wire_man_prod_w_lg_w_sum_one_range4232w5144w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5646w5652w5653w5654w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5646w5652w5653w(0) OR wire_man_prod_w_lg_w_sum_one_range4692w5650w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5657w5663w5664w5665w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5657w5663w5664w(0) OR wire_man_prod_w_lg_w_sum_one_range4702w5661w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5668w5674w5675w5676w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5668w5674w5675w(0) OR wire_man_prod_w_lg_w_sum_one_range4712w5672w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5679w5685w5686w5687w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5679w5685w5686w(0) OR wire_man_prod_w_lg_w_sum_one_range4722w5683w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5690w5696w5697w5698w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5690w5696w5697w(0) OR wire_man_prod_w_lg_w_sum_one_range4732w5694w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5701w5707w5708w5709w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5701w5707w5708w(0) OR wire_man_prod_w_lg_w_sum_one_range4742w5705w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5712w5718w5719w5720w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5712w5718w5719w(0) OR wire_man_prod_w_lg_w_sum_one_range4752w5716w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5723w5729w5730w5731w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5723w5729w5730w(0) OR wire_man_prod_w_lg_w_sum_one_range4762w5727w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5734w5740w5741w5742w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5734w5740w5741w(0) OR wire_man_prod_w_lg_w_sum_one_range4772w5738w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5745w5751w5752w5753w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5745w5751w5752w(0) OR wire_man_prod_w_lg_w_sum_one_range4782w5749w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5151w5157w5158w5159w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5151w5157w5158w(0) OR wire_man_prod_w_lg_w_sum_one_range4242w5155w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5756w5762w5763w5764w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5756w5762w5763w(0) OR wire_man_prod_w_lg_w_sum_one_range4792w5760w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5767w5773w5774w5775w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5767w5773w5774w(0) OR wire_man_prod_w_lg_w_sum_one_range4802w5771w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5778w5784w5785w5786w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5778w5784w5785w(0) OR wire_man_prod_w_lg_w_sum_one_range4812w5782w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5789w5795w5796w5797w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5789w5795w5796w(0) OR wire_man_prod_w_lg_w_sum_one_range4822w5793w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5800w5806w5807w5808w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5800w5806w5807w(0) OR wire_man_prod_w_lg_w_sum_one_range4832w5804w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5811w5817w5818w5819w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5811w5817w5818w(0) OR wire_man_prod_w_lg_w_sum_one_range4842w5815w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5822w5828w5829w5830w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5822w5828w5829w(0) OR wire_man_prod_w_lg_w_sum_one_range4852w5826w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5833w5839w5840w5841w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5833w5839w5840w(0) OR wire_man_prod_w_lg_w_sum_one_range4862w5837w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5844w5850w5851w5852w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5844w5850w5851w(0) OR wire_man_prod_w_lg_w_sum_one_range4872w5848w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5855w5861w5862w5863w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5855w5861w5862w(0) OR wire_man_prod_w_lg_w_sum_one_range4882w5859w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5162w5168w5169w5170w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5162w5168w5169w(0) OR wire_man_prod_w_lg_w_sum_one_range4252w5166w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5866w5872w5873w5874w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5866w5872w5873w(0) OR wire_man_prod_w_lg_w_sum_one_range4892w5870w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5877w5883w5884w5885w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5877w5883w5884w(0) OR wire_man_prod_w_lg_w_sum_one_range4902w5881w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5888w5894w5895w5896w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5888w5894w5895w(0) OR wire_man_prod_w_lg_w_sum_one_range4912w5892w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5899w5905w5906w5907w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5899w5905w5906w(0) OR wire_man_prod_w_lg_w_sum_one_range4922w5903w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5910w5916w5917w5918w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5910w5916w5917w(0) OR wire_man_prod_w_lg_w_sum_one_range4932w5914w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5921w5927w5928w5929w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5921w5927w5928w(0) OR wire_man_prod_w_lg_w_sum_one_range4942w5925w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5932w5938w5939w5940w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5932w5938w5939w(0) OR wire_man_prod_w_lg_w_sum_one_range4952w5936w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5943w5949w5950w5951w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5943w5949w5950w(0) OR wire_man_prod_w_lg_w_sum_one_range4962w5947w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5954w5960w5961w5962w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5954w5960w5961w(0) OR wire_man_prod_w_lg_w_sum_one_range4972w5958w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5965w5971w5972w5973w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5965w5971w5972w(0) OR wire_man_prod_w_lg_w_sum_one_range4982w5969w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5173w5179w5180w5181w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5173w5179w5180w(0) OR wire_man_prod_w_lg_w_sum_one_range4262w5177w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5976w5982w5983w5984w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5976w5982w5983w(0) OR wire_man_prod_w_lg_w_sum_one_range4992w5980w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5987w5993w5994w5995w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5987w5993w5994w(0) OR wire_man_prod_w_lg_w_sum_one_range5002w5991w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5998w6004w6005w6006w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5998w6004w6005w(0) OR wire_man_prod_w_lg_w_sum_one_range5012w6002w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6009w6015w6016w6017w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6009w6015w6016w(0) OR wire_man_prod_w_lg_w_sum_one_range5022w6013w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6020w6026w6027w6028w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6020w6026w6027w(0) OR wire_man_prod_w_lg_w_sum_one_range5032w6024w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6031w6037w6038w6039w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6031w6037w6038w(0) OR wire_man_prod_w_lg_w_sum_one_range5042w6035w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6042w6048w6049w6050w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6042w6048w6049w(0) OR wire_man_prod_w_lg_w_sum_one_range5052w6046w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6053w6059w6060w6061w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6053w6059w6060w(0) OR wire_man_prod_w_lg_w_sum_one_range5062w6057w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6064w6070w6071w6072w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6064w6070w6071w(0) OR wire_man_prod_w_lg_w_sum_one_range5072w6068w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6075w6081w6082w6083w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range6075w6081w6082w(0) OR wire_man_prod_w_lg_w_sum_one_range5082w6079w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5184w5190w5191w5192w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5184w5190w5191w(0) OR wire_man_prod_w_lg_w_sum_one_range4272w5188w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5195w5201w5202w5203w(0) <= wire_man_prod_w_lg_w_lg_w_vector1_range5195w5201w5202w(0) OR wire_man_prod_w_lg_w_sum_one_range4282w5199w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4187w4194w4195w4196w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4187w4194w4195w(0) OR wire_man_prod_w_lg_w_neg_msb_range4183w4192w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4289w4295w4296w4297w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4289w4295w4296w(0) OR wire_man_prod_w_lg_w_neg_msb_range4123w4293w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4299w4305w4306w4307w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4299w4305w4306w(0) OR wire_man_prod_w_lg_w_neg_msb_range4117w4303w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4309w4315w4316w4317w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4309w4315w4316w(0) OR wire_man_prod_w_lg_w_neg_msb_range4111w4313w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4319w4325w4326w4327w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4319w4325w4326w(0) OR wire_man_prod_w_lg_w_neg_msb_range4105w4323w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4329w4335w4336w4337w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4329w4335w4336w(0) OR wire_man_prod_w_lg_w_neg_msb_range4099w4333w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4339w4345w4346w4347w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4339w4345w4346w(0) OR wire_man_prod_w_lg_w_neg_msb_range4093w4343w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4349w4355w4356w4357w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4349w4355w4356w(0) OR wire_man_prod_w_lg_w_neg_msb_range4087w4353w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4359w4365w4366w4367w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4359w4365w4366w(0) OR wire_man_prod_w_lg_w_neg_msb_range4081w4363w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4369w4375w4376w4377w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4369w4375w4376w(0) OR wire_man_prod_w_lg_w_neg_msb_range4075w4373w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4379w4385w4386w4387w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4379w4385w4386w(0) OR wire_man_prod_w_lg_w_neg_msb_range4069w4383w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4199w4205w4206w4207w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4199w4205w4206w(0) OR wire_man_prod_w_lg_w_neg_msb_range4177w4203w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4389w4395w4396w4397w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4389w4395w4396w(0) OR wire_man_prod_w_lg_w_neg_msb_range4063w4393w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4399w4405w4406w4407w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4399w4405w4406w(0) OR wire_man_prod_w_lg_w_neg_msb_range4057w4403w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4409w4415w4416w4417w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4409w4415w4416w(0) OR wire_man_prod_w_lg_w_neg_msb_range4051w4413w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4419w4425w4426w4427w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4419w4425w4426w(0) OR wire_man_prod_w_lg_w_neg_msb_range4045w4423w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4429w4435w4436w4437w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4429w4435w4436w(0) OR wire_man_prod_w_lg_w_neg_msb_range4039w4433w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4439w4445w4446w4447w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4439w4445w4446w(0) OR wire_man_prod_w_lg_w_neg_msb_range4033w4443w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4449w4455w4456w4457w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4449w4455w4456w(0) OR wire_man_prod_w_lg_w_neg_msb_range4027w4453w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4459w4465w4466w4467w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4459w4465w4466w(0) OR wire_man_prod_w_lg_w_neg_msb_range4021w4463w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4469w4475w4476w4477w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4469w4475w4476w(0) OR wire_man_prod_w_lg_w_neg_msb_range4015w4473w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4479w4485w4486w4487w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4479w4485w4486w(0) OR wire_man_prod_w_lg_w_neg_msb_range4009w4483w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4209w4215w4216w4217w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4209w4215w4216w(0) OR wire_man_prod_w_lg_w_neg_msb_range4171w4213w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4489w4495w4496w4497w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4489w4495w4496w(0) OR wire_man_prod_w_lg_w_neg_msb_range4003w4493w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4499w4505w4506w4507w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4499w4505w4506w(0) OR wire_man_prod_w_lg_w_neg_msb_range3997w4503w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4509w4515w4516w4517w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4509w4515w4516w(0) OR wire_man_prod_w_lg_w_neg_msb_range3991w4513w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4519w4525w4526w4527w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4519w4525w4526w(0) OR wire_man_prod_w_lg_w_neg_msb_range3985w4523w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4529w4535w4536w4537w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4529w4535w4536w(0) OR wire_man_prod_w_lg_w_neg_msb_range3979w4533w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4539w4545w4546w4547w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4539w4545w4546w(0) OR wire_man_prod_w_lg_w_neg_msb_range3973w4543w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4549w4555w4556w4557w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4549w4555w4556w(0) OR wire_man_prod_w_lg_w_neg_msb_range3967w4553w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4559w4565w4566w4567w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4559w4565w4566w(0) OR wire_man_prod_w_lg_w_neg_msb_range3961w4563w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4569w4575w4576w4577w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4569w4575w4576w(0) OR wire_man_prod_w_lg_w_neg_msb_range3955w4573w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4579w4585w4586w4587w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4579w4585w4586w(0) OR wire_man_prod_w_lg_w_neg_msb_range3949w4583w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4219w4225w4226w4227w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4219w4225w4226w(0) OR wire_man_prod_w_lg_w_neg_msb_range4165w4223w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4589w4595w4596w4597w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4589w4595w4596w(0) OR wire_man_prod_w_lg_w_neg_msb_range3943w4593w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4599w4605w4606w4607w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4599w4605w4606w(0) OR wire_man_prod_w_lg_w_neg_msb_range3937w4603w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4609w4615w4616w4617w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4609w4615w4616w(0) OR wire_man_prod_w_lg_w_neg_msb_range3931w4613w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4619w4625w4626w4627w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4619w4625w4626w(0) OR wire_man_prod_w_lg_w_neg_msb_range3925w4623w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4629w4635w4636w4637w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4629w4635w4636w(0) OR wire_man_prod_w_lg_w_neg_msb_range3919w4633w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4639w4645w4646w4647w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4639w4645w4646w(0) OR wire_man_prod_w_lg_w_neg_msb_range3913w4643w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4649w4655w4656w4657w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4649w4655w4656w(0) OR wire_man_prod_w_lg_w_neg_msb_range3907w4653w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4659w4665w4666w4667w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4659w4665w4666w(0) OR wire_man_prod_w_lg_w_neg_msb_range3901w4663w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4669w4675w4676w4677w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4669w4675w4676w(0) OR wire_man_prod_w_lg_w_neg_msb_range3895w4673w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4679w4685w4686w4687w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4679w4685w4686w(0) OR wire_man_prod_w_lg_w_neg_msb_range3889w4683w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4229w4235w4236w4237w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4229w4235w4236w(0) OR wire_man_prod_w_lg_w_neg_msb_range4159w4233w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4689w4695w4696w4697w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4689w4695w4696w(0) OR wire_man_prod_w_lg_w_neg_msb_range3883w4693w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4699w4705w4706w4707w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4699w4705w4706w(0) OR wire_man_prod_w_lg_w_neg_msb_range3877w4703w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4709w4715w4716w4717w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4709w4715w4716w(0) OR wire_man_prod_w_lg_w_neg_msb_range3871w4713w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4719w4725w4726w4727w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4719w4725w4726w(0) OR wire_man_prod_w_lg_w_neg_msb_range3865w4723w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4729w4735w4736w4737w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4729w4735w4736w(0) OR wire_man_prod_w_lg_w_neg_msb_range3859w4733w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4739w4745w4746w4747w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4739w4745w4746w(0) OR wire_man_prod_w_lg_w_neg_msb_range3853w4743w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4749w4755w4756w4757w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4749w4755w4756w(0) OR wire_man_prod_w_lg_w_neg_msb_range3847w4753w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4759w4765w4766w4767w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4759w4765w4766w(0) OR wire_man_prod_w_lg_w_neg_msb_range3841w4763w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4769w4775w4776w4777w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4769w4775w4776w(0) OR wire_man_prod_w_lg_w_neg_msb_range3835w4773w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4779w4785w4786w4787w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4779w4785w4786w(0) OR wire_man_prod_w_lg_w_neg_msb_range3829w4783w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4239w4245w4246w4247w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4239w4245w4246w(0) OR wire_man_prod_w_lg_w_neg_msb_range4153w4243w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4789w4795w4796w4797w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4789w4795w4796w(0) OR wire_man_prod_w_lg_w_neg_msb_range3823w4793w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4799w4805w4806w4807w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4799w4805w4806w(0) OR wire_man_prod_w_lg_w_neg_msb_range3819w4803w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4809w4815w4816w4817w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4809w4815w4816w(0) OR wire_man_prod_w_lg_w_neg_msb_range3815w4813w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4819w4825w4826w4827w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4819w4825w4826w(0) OR wire_man_prod_w_lg_w_neg_msb_range3811w4823w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4829w4835w4836w4837w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4829w4835w4836w(0) OR wire_man_prod_w_lg_w_neg_msb_range3807w4833w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4839w4845w4846w4847w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4839w4845w4846w(0) OR wire_man_prod_w_lg_w_neg_msb_range3803w4843w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4849w4855w4856w4857w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4849w4855w4856w(0) OR wire_man_prod_w_lg_w_neg_msb_range3799w4853w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4859w4865w4866w4867w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4859w4865w4866w(0) OR wire_man_prod_w_lg_w_neg_msb_range3795w4863w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4869w4875w4876w4877w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4869w4875w4876w(0) OR wire_man_prod_w_lg_w_neg_msb_range3791w4873w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4879w4885w4886w4887w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4879w4885w4886w(0) OR wire_man_prod_w_lg_w_neg_msb_range3787w4883w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4249w4255w4256w4257w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4249w4255w4256w(0) OR wire_man_prod_w_lg_w_neg_msb_range4147w4253w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4889w4895w4896w4897w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4889w4895w4896w(0) OR wire_man_prod_w_lg_w_neg_msb_range3783w4893w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4899w4905w4906w4907w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4899w4905w4906w(0) OR wire_man_prod_w_lg_w_neg_msb_range3779w4903w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4909w4915w4916w4917w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4909w4915w4916w(0) OR wire_man_prod_w_lg_w_neg_msb_range3775w4913w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4919w4925w4926w4927w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4919w4925w4926w(0) OR wire_man_prod_w_lg_w_neg_msb_range3771w4923w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4929w4935w4936w4937w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4929w4935w4936w(0) OR wire_man_prod_w_lg_w_neg_msb_range3767w4933w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4939w4945w4946w4947w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4939w4945w4946w(0) OR wire_man_prod_w_lg_w_neg_msb_range3763w4943w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4949w4955w4956w4957w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4949w4955w4956w(0) OR wire_man_prod_w_lg_w_neg_msb_range3759w4953w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4959w4965w4966w4967w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4959w4965w4966w(0) OR wire_man_prod_w_lg_w_neg_msb_range3755w4963w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4969w4975w4976w4977w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4969w4975w4976w(0) OR wire_man_prod_w_lg_w_neg_msb_range3751w4973w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4979w4985w4986w4987w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4979w4985w4986w(0) OR wire_man_prod_w_lg_w_neg_msb_range3747w4983w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4259w4265w4266w4267w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4259w4265w4266w(0) OR wire_man_prod_w_lg_w_neg_msb_range4141w4263w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4989w4995w4996w4997w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4989w4995w4996w(0) OR wire_man_prod_w_lg_w_neg_msb_range3743w4993w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4999w5005w5006w5007w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4999w5005w5006w(0) OR wire_man_prod_w_lg_w_neg_msb_range3739w5003w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5009w5015w5016w5017w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5009w5015w5016w(0) OR wire_man_prod_w_lg_w_neg_msb_range3735w5013w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5019w5025w5026w5027w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5019w5025w5026w(0) OR wire_man_prod_w_lg_w_neg_msb_range3731w5023w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5029w5035w5036w5037w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5029w5035w5036w(0) OR wire_man_prod_w_lg_w_neg_msb_range3727w5033w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5039w5045w5046w5047w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5039w5045w5046w(0) OR wire_man_prod_w_lg_w_neg_msb_range3723w5043w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5049w5055w5056w5057w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5049w5055w5056w(0) OR wire_man_prod_w_lg_w_neg_msb_range3719w5053w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5059w5065w5066w5067w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5059w5065w5066w(0) OR wire_man_prod_w_lg_w_neg_msb_range3715w5063w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5069w5075w5076w5077w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5069w5075w5076w(0) OR wire_man_prod_w_lg_w_neg_msb_range3711w5073w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5079w5085w5086w5087w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range5079w5085w5086w(0) OR wire_man_prod_w_lg_w_neg_msb_range3705w5083w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4269w4275w4276w4277w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4269w4275w4276w(0) OR wire_man_prod_w_lg_w_neg_msb_range4135w4273w(0);
	wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4279w4285w4286w4287w(0) <= wire_man_prod_w_lg_w_lg_w_vector2_range4279w4285w4286w(0) OR wire_man_prod_w_lg_w_neg_msb_range4129w4283w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5094w5095w5096w(0) <= wire_man_prod_w_lg_w_vector1_range5094w5095w(0) XOR wire_man_prod_w_car_one_adj_range5092w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5206w5207w5208w(0) <= wire_man_prod_w_lg_w_vector1_range5206w5207w(0) XOR wire_man_prod_w_car_one_adj_range5205w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5217w5218w5219w(0) <= wire_man_prod_w_lg_w_vector1_range5217w5218w(0) XOR wire_man_prod_w_car_one_adj_range5216w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5228w5229w5230w(0) <= wire_man_prod_w_lg_w_vector1_range5228w5229w(0) XOR wire_man_prod_w_car_one_adj_range5227w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5239w5240w5241w(0) <= wire_man_prod_w_lg_w_vector1_range5239w5240w(0) XOR wire_man_prod_w_car_one_adj_range5238w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5250w5251w5252w(0) <= wire_man_prod_w_lg_w_vector1_range5250w5251w(0) XOR wire_man_prod_w_car_one_adj_range5249w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5261w5262w5263w(0) <= wire_man_prod_w_lg_w_vector1_range5261w5262w(0) XOR wire_man_prod_w_car_one_adj_range5260w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5272w5273w5274w(0) <= wire_man_prod_w_lg_w_vector1_range5272w5273w(0) XOR wire_man_prod_w_car_one_adj_range5271w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5283w5284w5285w(0) <= wire_man_prod_w_lg_w_vector1_range5283w5284w(0) XOR wire_man_prod_w_car_one_adj_range5282w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5294w5295w5296w(0) <= wire_man_prod_w_lg_w_vector1_range5294w5295w(0) XOR wire_man_prod_w_car_one_adj_range5293w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5305w5306w5307w(0) <= wire_man_prod_w_lg_w_vector1_range5305w5306w(0) XOR wire_man_prod_w_car_one_adj_range5304w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5107w5108w5109w(0) <= wire_man_prod_w_lg_w_vector1_range5107w5108w(0) XOR wire_man_prod_w_car_one_adj_range5106w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5316w5317w5318w(0) <= wire_man_prod_w_lg_w_vector1_range5316w5317w(0) XOR wire_man_prod_w_car_one_adj_range5315w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5327w5328w5329w(0) <= wire_man_prod_w_lg_w_vector1_range5327w5328w(0) XOR wire_man_prod_w_car_one_adj_range5326w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5338w5339w5340w(0) <= wire_man_prod_w_lg_w_vector1_range5338w5339w(0) XOR wire_man_prod_w_car_one_adj_range5337w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5349w5350w5351w(0) <= wire_man_prod_w_lg_w_vector1_range5349w5350w(0) XOR wire_man_prod_w_car_one_adj_range5348w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5360w5361w5362w(0) <= wire_man_prod_w_lg_w_vector1_range5360w5361w(0) XOR wire_man_prod_w_car_one_adj_range5359w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5371w5372w5373w(0) <= wire_man_prod_w_lg_w_vector1_range5371w5372w(0) XOR wire_man_prod_w_car_one_adj_range5370w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5382w5383w5384w(0) <= wire_man_prod_w_lg_w_vector1_range5382w5383w(0) XOR wire_man_prod_w_car_one_adj_range5381w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5393w5394w5395w(0) <= wire_man_prod_w_lg_w_vector1_range5393w5394w(0) XOR wire_man_prod_w_car_one_adj_range5392w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5404w5405w5406w(0) <= wire_man_prod_w_lg_w_vector1_range5404w5405w(0) XOR wire_man_prod_w_car_one_adj_range5403w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5415w5416w5417w(0) <= wire_man_prod_w_lg_w_vector1_range5415w5416w(0) XOR wire_man_prod_w_car_one_adj_range5414w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5118w5119w5120w(0) <= wire_man_prod_w_lg_w_vector1_range5118w5119w(0) XOR wire_man_prod_w_car_one_adj_range5117w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5426w5427w5428w(0) <= wire_man_prod_w_lg_w_vector1_range5426w5427w(0) XOR wire_man_prod_w_car_one_adj_range5425w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5437w5438w5439w(0) <= wire_man_prod_w_lg_w_vector1_range5437w5438w(0) XOR wire_man_prod_w_car_one_adj_range5436w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5448w5449w5450w(0) <= wire_man_prod_w_lg_w_vector1_range5448w5449w(0) XOR wire_man_prod_w_car_one_adj_range5447w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5459w5460w5461w(0) <= wire_man_prod_w_lg_w_vector1_range5459w5460w(0) XOR wire_man_prod_w_car_one_adj_range5458w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5470w5471w5472w(0) <= wire_man_prod_w_lg_w_vector1_range5470w5471w(0) XOR wire_man_prod_w_car_one_adj_range5469w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5481w5482w5483w(0) <= wire_man_prod_w_lg_w_vector1_range5481w5482w(0) XOR wire_man_prod_w_car_one_adj_range5480w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5492w5493w5494w(0) <= wire_man_prod_w_lg_w_vector1_range5492w5493w(0) XOR wire_man_prod_w_car_one_adj_range5491w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5503w5504w5505w(0) <= wire_man_prod_w_lg_w_vector1_range5503w5504w(0) XOR wire_man_prod_w_car_one_adj_range5502w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5514w5515w5516w(0) <= wire_man_prod_w_lg_w_vector1_range5514w5515w(0) XOR wire_man_prod_w_car_one_adj_range5513w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5525w5526w5527w(0) <= wire_man_prod_w_lg_w_vector1_range5525w5526w(0) XOR wire_man_prod_w_car_one_adj_range5524w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5129w5130w5131w(0) <= wire_man_prod_w_lg_w_vector1_range5129w5130w(0) XOR wire_man_prod_w_car_one_adj_range5128w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5536w5537w5538w(0) <= wire_man_prod_w_lg_w_vector1_range5536w5537w(0) XOR wire_man_prod_w_car_one_adj_range5535w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5547w5548w5549w(0) <= wire_man_prod_w_lg_w_vector1_range5547w5548w(0) XOR wire_man_prod_w_car_one_adj_range5546w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5558w5559w5560w(0) <= wire_man_prod_w_lg_w_vector1_range5558w5559w(0) XOR wire_man_prod_w_car_one_adj_range5557w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5569w5570w5571w(0) <= wire_man_prod_w_lg_w_vector1_range5569w5570w(0) XOR wire_man_prod_w_car_one_adj_range5568w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5580w5581w5582w(0) <= wire_man_prod_w_lg_w_vector1_range5580w5581w(0) XOR wire_man_prod_w_car_one_adj_range5579w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5591w5592w5593w(0) <= wire_man_prod_w_lg_w_vector1_range5591w5592w(0) XOR wire_man_prod_w_car_one_adj_range5590w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5602w5603w5604w(0) <= wire_man_prod_w_lg_w_vector1_range5602w5603w(0) XOR wire_man_prod_w_car_one_adj_range5601w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5613w5614w5615w(0) <= wire_man_prod_w_lg_w_vector1_range5613w5614w(0) XOR wire_man_prod_w_car_one_adj_range5612w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5624w5625w5626w(0) <= wire_man_prod_w_lg_w_vector1_range5624w5625w(0) XOR wire_man_prod_w_car_one_adj_range5623w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5635w5636w5637w(0) <= wire_man_prod_w_lg_w_vector1_range5635w5636w(0) XOR wire_man_prod_w_car_one_adj_range5634w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5140w5141w5142w(0) <= wire_man_prod_w_lg_w_vector1_range5140w5141w(0) XOR wire_man_prod_w_car_one_adj_range5139w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5646w5647w5648w(0) <= wire_man_prod_w_lg_w_vector1_range5646w5647w(0) XOR wire_man_prod_w_car_one_adj_range5645w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5657w5658w5659w(0) <= wire_man_prod_w_lg_w_vector1_range5657w5658w(0) XOR wire_man_prod_w_car_one_adj_range5656w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5668w5669w5670w(0) <= wire_man_prod_w_lg_w_vector1_range5668w5669w(0) XOR wire_man_prod_w_car_one_adj_range5667w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5679w5680w5681w(0) <= wire_man_prod_w_lg_w_vector1_range5679w5680w(0) XOR wire_man_prod_w_car_one_adj_range5678w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5690w5691w5692w(0) <= wire_man_prod_w_lg_w_vector1_range5690w5691w(0) XOR wire_man_prod_w_car_one_adj_range5689w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5701w5702w5703w(0) <= wire_man_prod_w_lg_w_vector1_range5701w5702w(0) XOR wire_man_prod_w_car_one_adj_range5700w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5712w5713w5714w(0) <= wire_man_prod_w_lg_w_vector1_range5712w5713w(0) XOR wire_man_prod_w_car_one_adj_range5711w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5723w5724w5725w(0) <= wire_man_prod_w_lg_w_vector1_range5723w5724w(0) XOR wire_man_prod_w_car_one_adj_range5722w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5734w5735w5736w(0) <= wire_man_prod_w_lg_w_vector1_range5734w5735w(0) XOR wire_man_prod_w_car_one_adj_range5733w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5745w5746w5747w(0) <= wire_man_prod_w_lg_w_vector1_range5745w5746w(0) XOR wire_man_prod_w_car_one_adj_range5744w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5151w5152w5153w(0) <= wire_man_prod_w_lg_w_vector1_range5151w5152w(0) XOR wire_man_prod_w_car_one_adj_range5150w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5756w5757w5758w(0) <= wire_man_prod_w_lg_w_vector1_range5756w5757w(0) XOR wire_man_prod_w_car_one_adj_range5755w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5767w5768w5769w(0) <= wire_man_prod_w_lg_w_vector1_range5767w5768w(0) XOR wire_man_prod_w_car_one_adj_range5766w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5778w5779w5780w(0) <= wire_man_prod_w_lg_w_vector1_range5778w5779w(0) XOR wire_man_prod_w_car_one_adj_range5777w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5789w5790w5791w(0) <= wire_man_prod_w_lg_w_vector1_range5789w5790w(0) XOR wire_man_prod_w_car_one_adj_range5788w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5800w5801w5802w(0) <= wire_man_prod_w_lg_w_vector1_range5800w5801w(0) XOR wire_man_prod_w_car_one_adj_range5799w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5811w5812w5813w(0) <= wire_man_prod_w_lg_w_vector1_range5811w5812w(0) XOR wire_man_prod_w_car_one_adj_range5810w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5822w5823w5824w(0) <= wire_man_prod_w_lg_w_vector1_range5822w5823w(0) XOR wire_man_prod_w_car_one_adj_range5821w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5833w5834w5835w(0) <= wire_man_prod_w_lg_w_vector1_range5833w5834w(0) XOR wire_man_prod_w_car_one_adj_range5832w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5844w5845w5846w(0) <= wire_man_prod_w_lg_w_vector1_range5844w5845w(0) XOR wire_man_prod_w_car_one_adj_range5843w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5855w5856w5857w(0) <= wire_man_prod_w_lg_w_vector1_range5855w5856w(0) XOR wire_man_prod_w_car_one_adj_range5854w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5162w5163w5164w(0) <= wire_man_prod_w_lg_w_vector1_range5162w5163w(0) XOR wire_man_prod_w_car_one_adj_range5161w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5866w5867w5868w(0) <= wire_man_prod_w_lg_w_vector1_range5866w5867w(0) XOR wire_man_prod_w_car_one_adj_range5865w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5877w5878w5879w(0) <= wire_man_prod_w_lg_w_vector1_range5877w5878w(0) XOR wire_man_prod_w_car_one_adj_range5876w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5888w5889w5890w(0) <= wire_man_prod_w_lg_w_vector1_range5888w5889w(0) XOR wire_man_prod_w_car_one_adj_range5887w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5899w5900w5901w(0) <= wire_man_prod_w_lg_w_vector1_range5899w5900w(0) XOR wire_man_prod_w_car_one_adj_range5898w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5910w5911w5912w(0) <= wire_man_prod_w_lg_w_vector1_range5910w5911w(0) XOR wire_man_prod_w_car_one_adj_range5909w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5921w5922w5923w(0) <= wire_man_prod_w_lg_w_vector1_range5921w5922w(0) XOR wire_man_prod_w_car_one_adj_range5920w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5932w5933w5934w(0) <= wire_man_prod_w_lg_w_vector1_range5932w5933w(0) XOR wire_man_prod_w_car_one_adj_range5931w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5943w5944w5945w(0) <= wire_man_prod_w_lg_w_vector1_range5943w5944w(0) XOR wire_man_prod_w_car_one_adj_range5942w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5954w5955w5956w(0) <= wire_man_prod_w_lg_w_vector1_range5954w5955w(0) XOR wire_man_prod_w_car_one_adj_range5953w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5965w5966w5967w(0) <= wire_man_prod_w_lg_w_vector1_range5965w5966w(0) XOR wire_man_prod_w_car_one_adj_range5964w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5173w5174w5175w(0) <= wire_man_prod_w_lg_w_vector1_range5173w5174w(0) XOR wire_man_prod_w_car_one_adj_range5172w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5976w5977w5978w(0) <= wire_man_prod_w_lg_w_vector1_range5976w5977w(0) XOR wire_man_prod_w_car_one_adj_range5975w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5987w5988w5989w(0) <= wire_man_prod_w_lg_w_vector1_range5987w5988w(0) XOR wire_man_prod_w_car_one_adj_range5986w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5998w5999w6000w(0) <= wire_man_prod_w_lg_w_vector1_range5998w5999w(0) XOR wire_man_prod_w_car_one_adj_range5997w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6009w6010w6011w(0) <= wire_man_prod_w_lg_w_vector1_range6009w6010w(0) XOR wire_man_prod_w_car_one_adj_range6008w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6020w6021w6022w(0) <= wire_man_prod_w_lg_w_vector1_range6020w6021w(0) XOR wire_man_prod_w_car_one_adj_range6019w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6031w6032w6033w(0) <= wire_man_prod_w_lg_w_vector1_range6031w6032w(0) XOR wire_man_prod_w_car_one_adj_range6030w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6042w6043w6044w(0) <= wire_man_prod_w_lg_w_vector1_range6042w6043w(0) XOR wire_man_prod_w_car_one_adj_range6041w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6053w6054w6055w(0) <= wire_man_prod_w_lg_w_vector1_range6053w6054w(0) XOR wire_man_prod_w_car_one_adj_range6052w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6064w6065w6066w(0) <= wire_man_prod_w_lg_w_vector1_range6064w6065w(0) XOR wire_man_prod_w_car_one_adj_range6063w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range6075w6076w6077w(0) <= wire_man_prod_w_lg_w_vector1_range6075w6076w(0) XOR wire_man_prod_w_car_one_adj_range6074w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5184w5185w5186w(0) <= wire_man_prod_w_lg_w_vector1_range5184w5185w(0) XOR wire_man_prod_w_car_one_adj_range5183w(0);
	wire_man_prod_w_lg_w_lg_w_vector1_range5195w5196w5197w(0) <= wire_man_prod_w_lg_w_vector1_range5195w5196w(0) XOR wire_man_prod_w_car_one_adj_range5194w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4187w4188w4189w(0) <= wire_man_prod_w_lg_w_vector2_range4187w4188w(0) XOR wire_man_prod_w_neg_lsb_range4186w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4289w4290w4291w(0) <= wire_man_prod_w_lg_w_vector2_range4289w4290w(0) XOR wire_man_prod_w_neg_lsb_range4126w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4299w4300w4301w(0) <= wire_man_prod_w_lg_w_vector2_range4299w4300w(0) XOR wire_man_prod_w_neg_lsb_range4120w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4309w4310w4311w(0) <= wire_man_prod_w_lg_w_vector2_range4309w4310w(0) XOR wire_man_prod_w_neg_lsb_range4114w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4319w4320w4321w(0) <= wire_man_prod_w_lg_w_vector2_range4319w4320w(0) XOR wire_man_prod_w_neg_lsb_range4108w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4329w4330w4331w(0) <= wire_man_prod_w_lg_w_vector2_range4329w4330w(0) XOR wire_man_prod_w_neg_lsb_range4102w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4339w4340w4341w(0) <= wire_man_prod_w_lg_w_vector2_range4339w4340w(0) XOR wire_man_prod_w_neg_lsb_range4096w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4349w4350w4351w(0) <= wire_man_prod_w_lg_w_vector2_range4349w4350w(0) XOR wire_man_prod_w_neg_lsb_range4090w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4359w4360w4361w(0) <= wire_man_prod_w_lg_w_vector2_range4359w4360w(0) XOR wire_man_prod_w_neg_lsb_range4084w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4369w4370w4371w(0) <= wire_man_prod_w_lg_w_vector2_range4369w4370w(0) XOR wire_man_prod_w_neg_lsb_range4078w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4379w4380w4381w(0) <= wire_man_prod_w_lg_w_vector2_range4379w4380w(0) XOR wire_man_prod_w_neg_lsb_range4072w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4199w4200w4201w(0) <= wire_man_prod_w_lg_w_vector2_range4199w4200w(0) XOR wire_man_prod_w_neg_lsb_range4180w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4389w4390w4391w(0) <= wire_man_prod_w_lg_w_vector2_range4389w4390w(0) XOR wire_man_prod_w_neg_lsb_range4066w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4399w4400w4401w(0) <= wire_man_prod_w_lg_w_vector2_range4399w4400w(0) XOR wire_man_prod_w_neg_lsb_range4060w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4409w4410w4411w(0) <= wire_man_prod_w_lg_w_vector2_range4409w4410w(0) XOR wire_man_prod_w_neg_lsb_range4054w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4419w4420w4421w(0) <= wire_man_prod_w_lg_w_vector2_range4419w4420w(0) XOR wire_man_prod_w_neg_lsb_range4048w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4429w4430w4431w(0) <= wire_man_prod_w_lg_w_vector2_range4429w4430w(0) XOR wire_man_prod_w_neg_lsb_range4042w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4439w4440w4441w(0) <= wire_man_prod_w_lg_w_vector2_range4439w4440w(0) XOR wire_man_prod_w_neg_lsb_range4036w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4449w4450w4451w(0) <= wire_man_prod_w_lg_w_vector2_range4449w4450w(0) XOR wire_man_prod_w_neg_lsb_range4030w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4459w4460w4461w(0) <= wire_man_prod_w_lg_w_vector2_range4459w4460w(0) XOR wire_man_prod_w_neg_lsb_range4024w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4469w4470w4471w(0) <= wire_man_prod_w_lg_w_vector2_range4469w4470w(0) XOR wire_man_prod_w_neg_lsb_range4018w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4479w4480w4481w(0) <= wire_man_prod_w_lg_w_vector2_range4479w4480w(0) XOR wire_man_prod_w_neg_lsb_range4012w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4209w4210w4211w(0) <= wire_man_prod_w_lg_w_vector2_range4209w4210w(0) XOR wire_man_prod_w_neg_lsb_range4174w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4489w4490w4491w(0) <= wire_man_prod_w_lg_w_vector2_range4489w4490w(0) XOR wire_man_prod_w_neg_lsb_range4006w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4499w4500w4501w(0) <= wire_man_prod_w_lg_w_vector2_range4499w4500w(0) XOR wire_man_prod_w_neg_lsb_range4000w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4509w4510w4511w(0) <= wire_man_prod_w_lg_w_vector2_range4509w4510w(0) XOR wire_man_prod_w_neg_lsb_range3994w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4519w4520w4521w(0) <= wire_man_prod_w_lg_w_vector2_range4519w4520w(0) XOR wire_man_prod_w_neg_lsb_range3988w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4529w4530w4531w(0) <= wire_man_prod_w_lg_w_vector2_range4529w4530w(0) XOR wire_man_prod_w_neg_lsb_range3982w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4539w4540w4541w(0) <= wire_man_prod_w_lg_w_vector2_range4539w4540w(0) XOR wire_man_prod_w_neg_lsb_range3976w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4549w4550w4551w(0) <= wire_man_prod_w_lg_w_vector2_range4549w4550w(0) XOR wire_man_prod_w_neg_lsb_range3970w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4559w4560w4561w(0) <= wire_man_prod_w_lg_w_vector2_range4559w4560w(0) XOR wire_man_prod_w_neg_lsb_range3964w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4569w4570w4571w(0) <= wire_man_prod_w_lg_w_vector2_range4569w4570w(0) XOR wire_man_prod_w_neg_lsb_range3958w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4579w4580w4581w(0) <= wire_man_prod_w_lg_w_vector2_range4579w4580w(0) XOR wire_man_prod_w_neg_lsb_range3952w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4219w4220w4221w(0) <= wire_man_prod_w_lg_w_vector2_range4219w4220w(0) XOR wire_man_prod_w_neg_lsb_range4168w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4589w4590w4591w(0) <= wire_man_prod_w_lg_w_vector2_range4589w4590w(0) XOR wire_man_prod_w_neg_lsb_range3946w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4599w4600w4601w(0) <= wire_man_prod_w_lg_w_vector2_range4599w4600w(0) XOR wire_man_prod_w_neg_lsb_range3940w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4609w4610w4611w(0) <= wire_man_prod_w_lg_w_vector2_range4609w4610w(0) XOR wire_man_prod_w_neg_lsb_range3934w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4619w4620w4621w(0) <= wire_man_prod_w_lg_w_vector2_range4619w4620w(0) XOR wire_man_prod_w_neg_lsb_range3928w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4629w4630w4631w(0) <= wire_man_prod_w_lg_w_vector2_range4629w4630w(0) XOR wire_man_prod_w_neg_lsb_range3922w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4639w4640w4641w(0) <= wire_man_prod_w_lg_w_vector2_range4639w4640w(0) XOR wire_man_prod_w_neg_lsb_range3916w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4649w4650w4651w(0) <= wire_man_prod_w_lg_w_vector2_range4649w4650w(0) XOR wire_man_prod_w_neg_lsb_range3910w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4659w4660w4661w(0) <= wire_man_prod_w_lg_w_vector2_range4659w4660w(0) XOR wire_man_prod_w_neg_lsb_range3904w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4669w4670w4671w(0) <= wire_man_prod_w_lg_w_vector2_range4669w4670w(0) XOR wire_man_prod_w_neg_lsb_range3898w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4679w4680w4681w(0) <= wire_man_prod_w_lg_w_vector2_range4679w4680w(0) XOR wire_man_prod_w_neg_lsb_range3892w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4229w4230w4231w(0) <= wire_man_prod_w_lg_w_vector2_range4229w4230w(0) XOR wire_man_prod_w_neg_lsb_range4162w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4689w4690w4691w(0) <= wire_man_prod_w_lg_w_vector2_range4689w4690w(0) XOR wire_man_prod_w_neg_lsb_range3886w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4699w4700w4701w(0) <= wire_man_prod_w_lg_w_vector2_range4699w4700w(0) XOR wire_man_prod_w_neg_lsb_range3880w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4709w4710w4711w(0) <= wire_man_prod_w_lg_w_vector2_range4709w4710w(0) XOR wire_man_prod_w_neg_lsb_range3874w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4719w4720w4721w(0) <= wire_man_prod_w_lg_w_vector2_range4719w4720w(0) XOR wire_man_prod_w_neg_lsb_range3868w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4729w4730w4731w(0) <= wire_man_prod_w_lg_w_vector2_range4729w4730w(0) XOR wire_man_prod_w_neg_lsb_range3862w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4739w4740w4741w(0) <= wire_man_prod_w_lg_w_vector2_range4739w4740w(0) XOR wire_man_prod_w_neg_lsb_range3856w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4749w4750w4751w(0) <= wire_man_prod_w_lg_w_vector2_range4749w4750w(0) XOR wire_man_prod_w_neg_lsb_range3850w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4759w4760w4761w(0) <= wire_man_prod_w_lg_w_vector2_range4759w4760w(0) XOR wire_man_prod_w_neg_lsb_range3844w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4769w4770w4771w(0) <= wire_man_prod_w_lg_w_vector2_range4769w4770w(0) XOR wire_man_prod_w_neg_lsb_range3838w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4779w4780w4781w(0) <= wire_man_prod_w_lg_w_vector2_range4779w4780w(0) XOR wire_man_prod_w_neg_lsb_range3832w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4239w4240w4241w(0) <= wire_man_prod_w_lg_w_vector2_range4239w4240w(0) XOR wire_man_prod_w_neg_lsb_range4156w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4789w4790w4791w(0) <= wire_man_prod_w_lg_w_vector2_range4789w4790w(0) XOR wire_man_prod_w_neg_lsb_range3825w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4799w4800w4801w(0) <= wire_man_prod_w_lg_w_vector2_range4799w4800w(0) XOR wire_man_prod_w_neg_lsb_range3821w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4809w4810w4811w(0) <= wire_man_prod_w_lg_w_vector2_range4809w4810w(0) XOR wire_man_prod_w_neg_lsb_range3817w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4819w4820w4821w(0) <= wire_man_prod_w_lg_w_vector2_range4819w4820w(0) XOR wire_man_prod_w_neg_lsb_range3813w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4829w4830w4831w(0) <= wire_man_prod_w_lg_w_vector2_range4829w4830w(0) XOR wire_man_prod_w_neg_lsb_range3809w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4839w4840w4841w(0) <= wire_man_prod_w_lg_w_vector2_range4839w4840w(0) XOR wire_man_prod_w_neg_lsb_range3805w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4849w4850w4851w(0) <= wire_man_prod_w_lg_w_vector2_range4849w4850w(0) XOR wire_man_prod_w_neg_lsb_range3801w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4859w4860w4861w(0) <= wire_man_prod_w_lg_w_vector2_range4859w4860w(0) XOR wire_man_prod_w_neg_lsb_range3797w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4869w4870w4871w(0) <= wire_man_prod_w_lg_w_vector2_range4869w4870w(0) XOR wire_man_prod_w_neg_lsb_range3793w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4879w4880w4881w(0) <= wire_man_prod_w_lg_w_vector2_range4879w4880w(0) XOR wire_man_prod_w_neg_lsb_range3789w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4249w4250w4251w(0) <= wire_man_prod_w_lg_w_vector2_range4249w4250w(0) XOR wire_man_prod_w_neg_lsb_range4150w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4889w4890w4891w(0) <= wire_man_prod_w_lg_w_vector2_range4889w4890w(0) XOR wire_man_prod_w_neg_lsb_range3785w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4899w4900w4901w(0) <= wire_man_prod_w_lg_w_vector2_range4899w4900w(0) XOR wire_man_prod_w_neg_lsb_range3781w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4909w4910w4911w(0) <= wire_man_prod_w_lg_w_vector2_range4909w4910w(0) XOR wire_man_prod_w_neg_lsb_range3777w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4919w4920w4921w(0) <= wire_man_prod_w_lg_w_vector2_range4919w4920w(0) XOR wire_man_prod_w_neg_lsb_range3773w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4929w4930w4931w(0) <= wire_man_prod_w_lg_w_vector2_range4929w4930w(0) XOR wire_man_prod_w_neg_lsb_range3769w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4939w4940w4941w(0) <= wire_man_prod_w_lg_w_vector2_range4939w4940w(0) XOR wire_man_prod_w_neg_lsb_range3765w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4949w4950w4951w(0) <= wire_man_prod_w_lg_w_vector2_range4949w4950w(0) XOR wire_man_prod_w_neg_lsb_range3761w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4959w4960w4961w(0) <= wire_man_prod_w_lg_w_vector2_range4959w4960w(0) XOR wire_man_prod_w_neg_lsb_range3757w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4969w4970w4971w(0) <= wire_man_prod_w_lg_w_vector2_range4969w4970w(0) XOR wire_man_prod_w_neg_lsb_range3753w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4979w4980w4981w(0) <= wire_man_prod_w_lg_w_vector2_range4979w4980w(0) XOR wire_man_prod_w_neg_lsb_range3749w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4259w4260w4261w(0) <= wire_man_prod_w_lg_w_vector2_range4259w4260w(0) XOR wire_man_prod_w_neg_lsb_range4144w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4989w4990w4991w(0) <= wire_man_prod_w_lg_w_vector2_range4989w4990w(0) XOR wire_man_prod_w_neg_lsb_range3745w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4999w5000w5001w(0) <= wire_man_prod_w_lg_w_vector2_range4999w5000w(0) XOR wire_man_prod_w_neg_lsb_range3741w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5009w5010w5011w(0) <= wire_man_prod_w_lg_w_vector2_range5009w5010w(0) XOR wire_man_prod_w_neg_lsb_range3737w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5019w5020w5021w(0) <= wire_man_prod_w_lg_w_vector2_range5019w5020w(0) XOR wire_man_prod_w_neg_lsb_range3733w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5029w5030w5031w(0) <= wire_man_prod_w_lg_w_vector2_range5029w5030w(0) XOR wire_man_prod_w_neg_lsb_range3729w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5039w5040w5041w(0) <= wire_man_prod_w_lg_w_vector2_range5039w5040w(0) XOR wire_man_prod_w_neg_lsb_range3725w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5049w5050w5051w(0) <= wire_man_prod_w_lg_w_vector2_range5049w5050w(0) XOR wire_man_prod_w_neg_lsb_range3721w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5059w5060w5061w(0) <= wire_man_prod_w_lg_w_vector2_range5059w5060w(0) XOR wire_man_prod_w_neg_lsb_range3717w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5069w5070w5071w(0) <= wire_man_prod_w_lg_w_vector2_range5069w5070w(0) XOR wire_man_prod_w_neg_lsb_range3713w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range5079w5080w5081w(0) <= wire_man_prod_w_lg_w_vector2_range5079w5080w(0) XOR wire_man_prod_w_neg_lsb_range3708w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4269w4270w4271w(0) <= wire_man_prod_w_lg_w_vector2_range4269w4270w(0) XOR wire_man_prod_w_neg_lsb_range4138w(0);
	wire_man_prod_w_lg_w_lg_w_vector2_range4279w4280w4281w(0) <= wire_man_prod_w_lg_w_vector2_range4279w4280w(0) XOR wire_man_prod_w_neg_lsb_range4132w(0);
	wire_man_prod_w_lg_w_vector1_range5094w5095w(0) <= wire_man_prod_w_vector1_range5094w(0) XOR wire_man_prod_w_sum_one_range4190w(0);
	wire_man_prod_w_lg_w_vector1_range5206w5207w(0) <= wire_man_prod_w_vector1_range5206w(0) XOR wire_man_prod_w_sum_one_range4292w(0);
	wire_man_prod_w_lg_w_vector1_range5217w5218w(0) <= wire_man_prod_w_vector1_range5217w(0) XOR wire_man_prod_w_sum_one_range4302w(0);
	wire_man_prod_w_lg_w_vector1_range5228w5229w(0) <= wire_man_prod_w_vector1_range5228w(0) XOR wire_man_prod_w_sum_one_range4312w(0);
	wire_man_prod_w_lg_w_vector1_range5239w5240w(0) <= wire_man_prod_w_vector1_range5239w(0) XOR wire_man_prod_w_sum_one_range4322w(0);
	wire_man_prod_w_lg_w_vector1_range5250w5251w(0) <= wire_man_prod_w_vector1_range5250w(0) XOR wire_man_prod_w_sum_one_range4332w(0);
	wire_man_prod_w_lg_w_vector1_range5261w5262w(0) <= wire_man_prod_w_vector1_range5261w(0) XOR wire_man_prod_w_sum_one_range4342w(0);
	wire_man_prod_w_lg_w_vector1_range5272w5273w(0) <= wire_man_prod_w_vector1_range5272w(0) XOR wire_man_prod_w_sum_one_range4352w(0);
	wire_man_prod_w_lg_w_vector1_range5283w5284w(0) <= wire_man_prod_w_vector1_range5283w(0) XOR wire_man_prod_w_sum_one_range4362w(0);
	wire_man_prod_w_lg_w_vector1_range5294w5295w(0) <= wire_man_prod_w_vector1_range5294w(0) XOR wire_man_prod_w_sum_one_range4372w(0);
	wire_man_prod_w_lg_w_vector1_range5305w5306w(0) <= wire_man_prod_w_vector1_range5305w(0) XOR wire_man_prod_w_sum_one_range4382w(0);
	wire_man_prod_w_lg_w_vector1_range5107w5108w(0) <= wire_man_prod_w_vector1_range5107w(0) XOR wire_man_prod_w_sum_one_range4202w(0);
	wire_man_prod_w_lg_w_vector1_range5316w5317w(0) <= wire_man_prod_w_vector1_range5316w(0) XOR wire_man_prod_w_sum_one_range4392w(0);
	wire_man_prod_w_lg_w_vector1_range5327w5328w(0) <= wire_man_prod_w_vector1_range5327w(0) XOR wire_man_prod_w_sum_one_range4402w(0);
	wire_man_prod_w_lg_w_vector1_range5338w5339w(0) <= wire_man_prod_w_vector1_range5338w(0) XOR wire_man_prod_w_sum_one_range4412w(0);
	wire_man_prod_w_lg_w_vector1_range5349w5350w(0) <= wire_man_prod_w_vector1_range5349w(0) XOR wire_man_prod_w_sum_one_range4422w(0);
	wire_man_prod_w_lg_w_vector1_range5360w5361w(0) <= wire_man_prod_w_vector1_range5360w(0) XOR wire_man_prod_w_sum_one_range4432w(0);
	wire_man_prod_w_lg_w_vector1_range5371w5372w(0) <= wire_man_prod_w_vector1_range5371w(0) XOR wire_man_prod_w_sum_one_range4442w(0);
	wire_man_prod_w_lg_w_vector1_range5382w5383w(0) <= wire_man_prod_w_vector1_range5382w(0) XOR wire_man_prod_w_sum_one_range4452w(0);
	wire_man_prod_w_lg_w_vector1_range5393w5394w(0) <= wire_man_prod_w_vector1_range5393w(0) XOR wire_man_prod_w_sum_one_range4462w(0);
	wire_man_prod_w_lg_w_vector1_range5404w5405w(0) <= wire_man_prod_w_vector1_range5404w(0) XOR wire_man_prod_w_sum_one_range4472w(0);
	wire_man_prod_w_lg_w_vector1_range5415w5416w(0) <= wire_man_prod_w_vector1_range5415w(0) XOR wire_man_prod_w_sum_one_range4482w(0);
	wire_man_prod_w_lg_w_vector1_range5118w5119w(0) <= wire_man_prod_w_vector1_range5118w(0) XOR wire_man_prod_w_sum_one_range4212w(0);
	wire_man_prod_w_lg_w_vector1_range5426w5427w(0) <= wire_man_prod_w_vector1_range5426w(0) XOR wire_man_prod_w_sum_one_range4492w(0);
	wire_man_prod_w_lg_w_vector1_range5437w5438w(0) <= wire_man_prod_w_vector1_range5437w(0) XOR wire_man_prod_w_sum_one_range4502w(0);
	wire_man_prod_w_lg_w_vector1_range5448w5449w(0) <= wire_man_prod_w_vector1_range5448w(0) XOR wire_man_prod_w_sum_one_range4512w(0);
	wire_man_prod_w_lg_w_vector1_range5459w5460w(0) <= wire_man_prod_w_vector1_range5459w(0) XOR wire_man_prod_w_sum_one_range4522w(0);
	wire_man_prod_w_lg_w_vector1_range5470w5471w(0) <= wire_man_prod_w_vector1_range5470w(0) XOR wire_man_prod_w_sum_one_range4532w(0);
	wire_man_prod_w_lg_w_vector1_range5481w5482w(0) <= wire_man_prod_w_vector1_range5481w(0) XOR wire_man_prod_w_sum_one_range4542w(0);
	wire_man_prod_w_lg_w_vector1_range5492w5493w(0) <= wire_man_prod_w_vector1_range5492w(0) XOR wire_man_prod_w_sum_one_range4552w(0);
	wire_man_prod_w_lg_w_vector1_range5503w5504w(0) <= wire_man_prod_w_vector1_range5503w(0) XOR wire_man_prod_w_sum_one_range4562w(0);
	wire_man_prod_w_lg_w_vector1_range5514w5515w(0) <= wire_man_prod_w_vector1_range5514w(0) XOR wire_man_prod_w_sum_one_range4572w(0);
	wire_man_prod_w_lg_w_vector1_range5525w5526w(0) <= wire_man_prod_w_vector1_range5525w(0) XOR wire_man_prod_w_sum_one_range4582w(0);
	wire_man_prod_w_lg_w_vector1_range5129w5130w(0) <= wire_man_prod_w_vector1_range5129w(0) XOR wire_man_prod_w_sum_one_range4222w(0);
	wire_man_prod_w_lg_w_vector1_range5536w5537w(0) <= wire_man_prod_w_vector1_range5536w(0) XOR wire_man_prod_w_sum_one_range4592w(0);
	wire_man_prod_w_lg_w_vector1_range5547w5548w(0) <= wire_man_prod_w_vector1_range5547w(0) XOR wire_man_prod_w_sum_one_range4602w(0);
	wire_man_prod_w_lg_w_vector1_range5558w5559w(0) <= wire_man_prod_w_vector1_range5558w(0) XOR wire_man_prod_w_sum_one_range4612w(0);
	wire_man_prod_w_lg_w_vector1_range5569w5570w(0) <= wire_man_prod_w_vector1_range5569w(0) XOR wire_man_prod_w_sum_one_range4622w(0);
	wire_man_prod_w_lg_w_vector1_range5580w5581w(0) <= wire_man_prod_w_vector1_range5580w(0) XOR wire_man_prod_w_sum_one_range4632w(0);
	wire_man_prod_w_lg_w_vector1_range5591w5592w(0) <= wire_man_prod_w_vector1_range5591w(0) XOR wire_man_prod_w_sum_one_range4642w(0);
	wire_man_prod_w_lg_w_vector1_range5602w5603w(0) <= wire_man_prod_w_vector1_range5602w(0) XOR wire_man_prod_w_sum_one_range4652w(0);
	wire_man_prod_w_lg_w_vector1_range5613w5614w(0) <= wire_man_prod_w_vector1_range5613w(0) XOR wire_man_prod_w_sum_one_range4662w(0);
	wire_man_prod_w_lg_w_vector1_range5624w5625w(0) <= wire_man_prod_w_vector1_range5624w(0) XOR wire_man_prod_w_sum_one_range4672w(0);
	wire_man_prod_w_lg_w_vector1_range5635w5636w(0) <= wire_man_prod_w_vector1_range5635w(0) XOR wire_man_prod_w_sum_one_range4682w(0);
	wire_man_prod_w_lg_w_vector1_range5140w5141w(0) <= wire_man_prod_w_vector1_range5140w(0) XOR wire_man_prod_w_sum_one_range4232w(0);
	wire_man_prod_w_lg_w_vector1_range5646w5647w(0) <= wire_man_prod_w_vector1_range5646w(0) XOR wire_man_prod_w_sum_one_range4692w(0);
	wire_man_prod_w_lg_w_vector1_range5657w5658w(0) <= wire_man_prod_w_vector1_range5657w(0) XOR wire_man_prod_w_sum_one_range4702w(0);
	wire_man_prod_w_lg_w_vector1_range5668w5669w(0) <= wire_man_prod_w_vector1_range5668w(0) XOR wire_man_prod_w_sum_one_range4712w(0);
	wire_man_prod_w_lg_w_vector1_range5679w5680w(0) <= wire_man_prod_w_vector1_range5679w(0) XOR wire_man_prod_w_sum_one_range4722w(0);
	wire_man_prod_w_lg_w_vector1_range5690w5691w(0) <= wire_man_prod_w_vector1_range5690w(0) XOR wire_man_prod_w_sum_one_range4732w(0);
	wire_man_prod_w_lg_w_vector1_range5701w5702w(0) <= wire_man_prod_w_vector1_range5701w(0) XOR wire_man_prod_w_sum_one_range4742w(0);
	wire_man_prod_w_lg_w_vector1_range5712w5713w(0) <= wire_man_prod_w_vector1_range5712w(0) XOR wire_man_prod_w_sum_one_range4752w(0);
	wire_man_prod_w_lg_w_vector1_range5723w5724w(0) <= wire_man_prod_w_vector1_range5723w(0) XOR wire_man_prod_w_sum_one_range4762w(0);
	wire_man_prod_w_lg_w_vector1_range5734w5735w(0) <= wire_man_prod_w_vector1_range5734w(0) XOR wire_man_prod_w_sum_one_range4772w(0);
	wire_man_prod_w_lg_w_vector1_range5745w5746w(0) <= wire_man_prod_w_vector1_range5745w(0) XOR wire_man_prod_w_sum_one_range4782w(0);
	wire_man_prod_w_lg_w_vector1_range5151w5152w(0) <= wire_man_prod_w_vector1_range5151w(0) XOR wire_man_prod_w_sum_one_range4242w(0);
	wire_man_prod_w_lg_w_vector1_range5756w5757w(0) <= wire_man_prod_w_vector1_range5756w(0) XOR wire_man_prod_w_sum_one_range4792w(0);
	wire_man_prod_w_lg_w_vector1_range5767w5768w(0) <= wire_man_prod_w_vector1_range5767w(0) XOR wire_man_prod_w_sum_one_range4802w(0);
	wire_man_prod_w_lg_w_vector1_range5778w5779w(0) <= wire_man_prod_w_vector1_range5778w(0) XOR wire_man_prod_w_sum_one_range4812w(0);
	wire_man_prod_w_lg_w_vector1_range5789w5790w(0) <= wire_man_prod_w_vector1_range5789w(0) XOR wire_man_prod_w_sum_one_range4822w(0);
	wire_man_prod_w_lg_w_vector1_range5800w5801w(0) <= wire_man_prod_w_vector1_range5800w(0) XOR wire_man_prod_w_sum_one_range4832w(0);
	wire_man_prod_w_lg_w_vector1_range5811w5812w(0) <= wire_man_prod_w_vector1_range5811w(0) XOR wire_man_prod_w_sum_one_range4842w(0);
	wire_man_prod_w_lg_w_vector1_range5822w5823w(0) <= wire_man_prod_w_vector1_range5822w(0) XOR wire_man_prod_w_sum_one_range4852w(0);
	wire_man_prod_w_lg_w_vector1_range5833w5834w(0) <= wire_man_prod_w_vector1_range5833w(0) XOR wire_man_prod_w_sum_one_range4862w(0);
	wire_man_prod_w_lg_w_vector1_range5844w5845w(0) <= wire_man_prod_w_vector1_range5844w(0) XOR wire_man_prod_w_sum_one_range4872w(0);
	wire_man_prod_w_lg_w_vector1_range5855w5856w(0) <= wire_man_prod_w_vector1_range5855w(0) XOR wire_man_prod_w_sum_one_range4882w(0);
	wire_man_prod_w_lg_w_vector1_range5162w5163w(0) <= wire_man_prod_w_vector1_range5162w(0) XOR wire_man_prod_w_sum_one_range4252w(0);
	wire_man_prod_w_lg_w_vector1_range5866w5867w(0) <= wire_man_prod_w_vector1_range5866w(0) XOR wire_man_prod_w_sum_one_range4892w(0);
	wire_man_prod_w_lg_w_vector1_range5877w5878w(0) <= wire_man_prod_w_vector1_range5877w(0) XOR wire_man_prod_w_sum_one_range4902w(0);
	wire_man_prod_w_lg_w_vector1_range5888w5889w(0) <= wire_man_prod_w_vector1_range5888w(0) XOR wire_man_prod_w_sum_one_range4912w(0);
	wire_man_prod_w_lg_w_vector1_range5899w5900w(0) <= wire_man_prod_w_vector1_range5899w(0) XOR wire_man_prod_w_sum_one_range4922w(0);
	wire_man_prod_w_lg_w_vector1_range5910w5911w(0) <= wire_man_prod_w_vector1_range5910w(0) XOR wire_man_prod_w_sum_one_range4932w(0);
	wire_man_prod_w_lg_w_vector1_range5921w5922w(0) <= wire_man_prod_w_vector1_range5921w(0) XOR wire_man_prod_w_sum_one_range4942w(0);
	wire_man_prod_w_lg_w_vector1_range5932w5933w(0) <= wire_man_prod_w_vector1_range5932w(0) XOR wire_man_prod_w_sum_one_range4952w(0);
	wire_man_prod_w_lg_w_vector1_range5943w5944w(0) <= wire_man_prod_w_vector1_range5943w(0) XOR wire_man_prod_w_sum_one_range4962w(0);
	wire_man_prod_w_lg_w_vector1_range5954w5955w(0) <= wire_man_prod_w_vector1_range5954w(0) XOR wire_man_prod_w_sum_one_range4972w(0);
	wire_man_prod_w_lg_w_vector1_range5965w5966w(0) <= wire_man_prod_w_vector1_range5965w(0) XOR wire_man_prod_w_sum_one_range4982w(0);
	wire_man_prod_w_lg_w_vector1_range5173w5174w(0) <= wire_man_prod_w_vector1_range5173w(0) XOR wire_man_prod_w_sum_one_range4262w(0);
	wire_man_prod_w_lg_w_vector1_range5976w5977w(0) <= wire_man_prod_w_vector1_range5976w(0) XOR wire_man_prod_w_sum_one_range4992w(0);
	wire_man_prod_w_lg_w_vector1_range5987w5988w(0) <= wire_man_prod_w_vector1_range5987w(0) XOR wire_man_prod_w_sum_one_range5002w(0);
	wire_man_prod_w_lg_w_vector1_range5998w5999w(0) <= wire_man_prod_w_vector1_range5998w(0) XOR wire_man_prod_w_sum_one_range5012w(0);
	wire_man_prod_w_lg_w_vector1_range6009w6010w(0) <= wire_man_prod_w_vector1_range6009w(0) XOR wire_man_prod_w_sum_one_range5022w(0);
	wire_man_prod_w_lg_w_vector1_range6020w6021w(0) <= wire_man_prod_w_vector1_range6020w(0) XOR wire_man_prod_w_sum_one_range5032w(0);
	wire_man_prod_w_lg_w_vector1_range6031w6032w(0) <= wire_man_prod_w_vector1_range6031w(0) XOR wire_man_prod_w_sum_one_range5042w(0);
	wire_man_prod_w_lg_w_vector1_range6042w6043w(0) <= wire_man_prod_w_vector1_range6042w(0) XOR wire_man_prod_w_sum_one_range5052w(0);
	wire_man_prod_w_lg_w_vector1_range6053w6054w(0) <= wire_man_prod_w_vector1_range6053w(0) XOR wire_man_prod_w_sum_one_range5062w(0);
	wire_man_prod_w_lg_w_vector1_range6064w6065w(0) <= wire_man_prod_w_vector1_range6064w(0) XOR wire_man_prod_w_sum_one_range5072w(0);
	wire_man_prod_w_lg_w_vector1_range6075w6076w(0) <= wire_man_prod_w_vector1_range6075w(0) XOR wire_man_prod_w_sum_one_range5082w(0);
	wire_man_prod_w_lg_w_vector1_range5184w5185w(0) <= wire_man_prod_w_vector1_range5184w(0) XOR wire_man_prod_w_sum_one_range4272w(0);
	wire_man_prod_w_lg_w_vector1_range5195w5196w(0) <= wire_man_prod_w_vector1_range5195w(0) XOR wire_man_prod_w_sum_one_range4282w(0);
	wire_man_prod_w_lg_w_vector2_range4187w4188w(0) <= wire_man_prod_w_vector2_range4187w(0) XOR wire_man_prod_w_neg_msb_range4183w(0);
	wire_man_prod_w_lg_w_vector2_range4289w4290w(0) <= wire_man_prod_w_vector2_range4289w(0) XOR wire_man_prod_w_neg_msb_range4123w(0);
	wire_man_prod_w_lg_w_vector2_range4299w4300w(0) <= wire_man_prod_w_vector2_range4299w(0) XOR wire_man_prod_w_neg_msb_range4117w(0);
	wire_man_prod_w_lg_w_vector2_range4309w4310w(0) <= wire_man_prod_w_vector2_range4309w(0) XOR wire_man_prod_w_neg_msb_range4111w(0);
	wire_man_prod_w_lg_w_vector2_range4319w4320w(0) <= wire_man_prod_w_vector2_range4319w(0) XOR wire_man_prod_w_neg_msb_range4105w(0);
	wire_man_prod_w_lg_w_vector2_range4329w4330w(0) <= wire_man_prod_w_vector2_range4329w(0) XOR wire_man_prod_w_neg_msb_range4099w(0);
	wire_man_prod_w_lg_w_vector2_range4339w4340w(0) <= wire_man_prod_w_vector2_range4339w(0) XOR wire_man_prod_w_neg_msb_range4093w(0);
	wire_man_prod_w_lg_w_vector2_range4349w4350w(0) <= wire_man_prod_w_vector2_range4349w(0) XOR wire_man_prod_w_neg_msb_range4087w(0);
	wire_man_prod_w_lg_w_vector2_range4359w4360w(0) <= wire_man_prod_w_vector2_range4359w(0) XOR wire_man_prod_w_neg_msb_range4081w(0);
	wire_man_prod_w_lg_w_vector2_range4369w4370w(0) <= wire_man_prod_w_vector2_range4369w(0) XOR wire_man_prod_w_neg_msb_range4075w(0);
	wire_man_prod_w_lg_w_vector2_range4379w4380w(0) <= wire_man_prod_w_vector2_range4379w(0) XOR wire_man_prod_w_neg_msb_range4069w(0);
	wire_man_prod_w_lg_w_vector2_range4199w4200w(0) <= wire_man_prod_w_vector2_range4199w(0) XOR wire_man_prod_w_neg_msb_range4177w(0);
	wire_man_prod_w_lg_w_vector2_range4389w4390w(0) <= wire_man_prod_w_vector2_range4389w(0) XOR wire_man_prod_w_neg_msb_range4063w(0);
	wire_man_prod_w_lg_w_vector2_range4399w4400w(0) <= wire_man_prod_w_vector2_range4399w(0) XOR wire_man_prod_w_neg_msb_range4057w(0);
	wire_man_prod_w_lg_w_vector2_range4409w4410w(0) <= wire_man_prod_w_vector2_range4409w(0) XOR wire_man_prod_w_neg_msb_range4051w(0);
	wire_man_prod_w_lg_w_vector2_range4419w4420w(0) <= wire_man_prod_w_vector2_range4419w(0) XOR wire_man_prod_w_neg_msb_range4045w(0);
	wire_man_prod_w_lg_w_vector2_range4429w4430w(0) <= wire_man_prod_w_vector2_range4429w(0) XOR wire_man_prod_w_neg_msb_range4039w(0);
	wire_man_prod_w_lg_w_vector2_range4439w4440w(0) <= wire_man_prod_w_vector2_range4439w(0) XOR wire_man_prod_w_neg_msb_range4033w(0);
	wire_man_prod_w_lg_w_vector2_range4449w4450w(0) <= wire_man_prod_w_vector2_range4449w(0) XOR wire_man_prod_w_neg_msb_range4027w(0);
	wire_man_prod_w_lg_w_vector2_range4459w4460w(0) <= wire_man_prod_w_vector2_range4459w(0) XOR wire_man_prod_w_neg_msb_range4021w(0);
	wire_man_prod_w_lg_w_vector2_range4469w4470w(0) <= wire_man_prod_w_vector2_range4469w(0) XOR wire_man_prod_w_neg_msb_range4015w(0);
	wire_man_prod_w_lg_w_vector2_range4479w4480w(0) <= wire_man_prod_w_vector2_range4479w(0) XOR wire_man_prod_w_neg_msb_range4009w(0);
	wire_man_prod_w_lg_w_vector2_range4209w4210w(0) <= wire_man_prod_w_vector2_range4209w(0) XOR wire_man_prod_w_neg_msb_range4171w(0);
	wire_man_prod_w_lg_w_vector2_range4489w4490w(0) <= wire_man_prod_w_vector2_range4489w(0) XOR wire_man_prod_w_neg_msb_range4003w(0);
	wire_man_prod_w_lg_w_vector2_range4499w4500w(0) <= wire_man_prod_w_vector2_range4499w(0) XOR wire_man_prod_w_neg_msb_range3997w(0);
	wire_man_prod_w_lg_w_vector2_range4509w4510w(0) <= wire_man_prod_w_vector2_range4509w(0) XOR wire_man_prod_w_neg_msb_range3991w(0);
	wire_man_prod_w_lg_w_vector2_range4519w4520w(0) <= wire_man_prod_w_vector2_range4519w(0) XOR wire_man_prod_w_neg_msb_range3985w(0);
	wire_man_prod_w_lg_w_vector2_range4529w4530w(0) <= wire_man_prod_w_vector2_range4529w(0) XOR wire_man_prod_w_neg_msb_range3979w(0);
	wire_man_prod_w_lg_w_vector2_range4539w4540w(0) <= wire_man_prod_w_vector2_range4539w(0) XOR wire_man_prod_w_neg_msb_range3973w(0);
	wire_man_prod_w_lg_w_vector2_range4549w4550w(0) <= wire_man_prod_w_vector2_range4549w(0) XOR wire_man_prod_w_neg_msb_range3967w(0);
	wire_man_prod_w_lg_w_vector2_range4559w4560w(0) <= wire_man_prod_w_vector2_range4559w(0) XOR wire_man_prod_w_neg_msb_range3961w(0);
	wire_man_prod_w_lg_w_vector2_range4569w4570w(0) <= wire_man_prod_w_vector2_range4569w(0) XOR wire_man_prod_w_neg_msb_range3955w(0);
	wire_man_prod_w_lg_w_vector2_range4579w4580w(0) <= wire_man_prod_w_vector2_range4579w(0) XOR wire_man_prod_w_neg_msb_range3949w(0);
	wire_man_prod_w_lg_w_vector2_range4219w4220w(0) <= wire_man_prod_w_vector2_range4219w(0) XOR wire_man_prod_w_neg_msb_range4165w(0);
	wire_man_prod_w_lg_w_vector2_range4589w4590w(0) <= wire_man_prod_w_vector2_range4589w(0) XOR wire_man_prod_w_neg_msb_range3943w(0);
	wire_man_prod_w_lg_w_vector2_range4599w4600w(0) <= wire_man_prod_w_vector2_range4599w(0) XOR wire_man_prod_w_neg_msb_range3937w(0);
	wire_man_prod_w_lg_w_vector2_range4609w4610w(0) <= wire_man_prod_w_vector2_range4609w(0) XOR wire_man_prod_w_neg_msb_range3931w(0);
	wire_man_prod_w_lg_w_vector2_range4619w4620w(0) <= wire_man_prod_w_vector2_range4619w(0) XOR wire_man_prod_w_neg_msb_range3925w(0);
	wire_man_prod_w_lg_w_vector2_range4629w4630w(0) <= wire_man_prod_w_vector2_range4629w(0) XOR wire_man_prod_w_neg_msb_range3919w(0);
	wire_man_prod_w_lg_w_vector2_range4639w4640w(0) <= wire_man_prod_w_vector2_range4639w(0) XOR wire_man_prod_w_neg_msb_range3913w(0);
	wire_man_prod_w_lg_w_vector2_range4649w4650w(0) <= wire_man_prod_w_vector2_range4649w(0) XOR wire_man_prod_w_neg_msb_range3907w(0);
	wire_man_prod_w_lg_w_vector2_range4659w4660w(0) <= wire_man_prod_w_vector2_range4659w(0) XOR wire_man_prod_w_neg_msb_range3901w(0);
	wire_man_prod_w_lg_w_vector2_range4669w4670w(0) <= wire_man_prod_w_vector2_range4669w(0) XOR wire_man_prod_w_neg_msb_range3895w(0);
	wire_man_prod_w_lg_w_vector2_range4679w4680w(0) <= wire_man_prod_w_vector2_range4679w(0) XOR wire_man_prod_w_neg_msb_range3889w(0);
	wire_man_prod_w_lg_w_vector2_range4229w4230w(0) <= wire_man_prod_w_vector2_range4229w(0) XOR wire_man_prod_w_neg_msb_range4159w(0);
	wire_man_prod_w_lg_w_vector2_range4689w4690w(0) <= wire_man_prod_w_vector2_range4689w(0) XOR wire_man_prod_w_neg_msb_range3883w(0);
	wire_man_prod_w_lg_w_vector2_range4699w4700w(0) <= wire_man_prod_w_vector2_range4699w(0) XOR wire_man_prod_w_neg_msb_range3877w(0);
	wire_man_prod_w_lg_w_vector2_range4709w4710w(0) <= wire_man_prod_w_vector2_range4709w(0) XOR wire_man_prod_w_neg_msb_range3871w(0);
	wire_man_prod_w_lg_w_vector2_range4719w4720w(0) <= wire_man_prod_w_vector2_range4719w(0) XOR wire_man_prod_w_neg_msb_range3865w(0);
	wire_man_prod_w_lg_w_vector2_range4729w4730w(0) <= wire_man_prod_w_vector2_range4729w(0) XOR wire_man_prod_w_neg_msb_range3859w(0);
	wire_man_prod_w_lg_w_vector2_range4739w4740w(0) <= wire_man_prod_w_vector2_range4739w(0) XOR wire_man_prod_w_neg_msb_range3853w(0);
	wire_man_prod_w_lg_w_vector2_range4749w4750w(0) <= wire_man_prod_w_vector2_range4749w(0) XOR wire_man_prod_w_neg_msb_range3847w(0);
	wire_man_prod_w_lg_w_vector2_range4759w4760w(0) <= wire_man_prod_w_vector2_range4759w(0) XOR wire_man_prod_w_neg_msb_range3841w(0);
	wire_man_prod_w_lg_w_vector2_range4769w4770w(0) <= wire_man_prod_w_vector2_range4769w(0) XOR wire_man_prod_w_neg_msb_range3835w(0);
	wire_man_prod_w_lg_w_vector2_range4779w4780w(0) <= wire_man_prod_w_vector2_range4779w(0) XOR wire_man_prod_w_neg_msb_range3829w(0);
	wire_man_prod_w_lg_w_vector2_range4239w4240w(0) <= wire_man_prod_w_vector2_range4239w(0) XOR wire_man_prod_w_neg_msb_range4153w(0);
	wire_man_prod_w_lg_w_vector2_range4789w4790w(0) <= wire_man_prod_w_vector2_range4789w(0) XOR wire_man_prod_w_neg_msb_range3823w(0);
	wire_man_prod_w_lg_w_vector2_range4799w4800w(0) <= wire_man_prod_w_vector2_range4799w(0) XOR wire_man_prod_w_neg_msb_range3819w(0);
	wire_man_prod_w_lg_w_vector2_range4809w4810w(0) <= wire_man_prod_w_vector2_range4809w(0) XOR wire_man_prod_w_neg_msb_range3815w(0);
	wire_man_prod_w_lg_w_vector2_range4819w4820w(0) <= wire_man_prod_w_vector2_range4819w(0) XOR wire_man_prod_w_neg_msb_range3811w(0);
	wire_man_prod_w_lg_w_vector2_range4829w4830w(0) <= wire_man_prod_w_vector2_range4829w(0) XOR wire_man_prod_w_neg_msb_range3807w(0);
	wire_man_prod_w_lg_w_vector2_range4839w4840w(0) <= wire_man_prod_w_vector2_range4839w(0) XOR wire_man_prod_w_neg_msb_range3803w(0);
	wire_man_prod_w_lg_w_vector2_range4849w4850w(0) <= wire_man_prod_w_vector2_range4849w(0) XOR wire_man_prod_w_neg_msb_range3799w(0);
	wire_man_prod_w_lg_w_vector2_range4859w4860w(0) <= wire_man_prod_w_vector2_range4859w(0) XOR wire_man_prod_w_neg_msb_range3795w(0);
	wire_man_prod_w_lg_w_vector2_range4869w4870w(0) <= wire_man_prod_w_vector2_range4869w(0) XOR wire_man_prod_w_neg_msb_range3791w(0);
	wire_man_prod_w_lg_w_vector2_range4879w4880w(0) <= wire_man_prod_w_vector2_range4879w(0) XOR wire_man_prod_w_neg_msb_range3787w(0);
	wire_man_prod_w_lg_w_vector2_range4249w4250w(0) <= wire_man_prod_w_vector2_range4249w(0) XOR wire_man_prod_w_neg_msb_range4147w(0);
	wire_man_prod_w_lg_w_vector2_range4889w4890w(0) <= wire_man_prod_w_vector2_range4889w(0) XOR wire_man_prod_w_neg_msb_range3783w(0);
	wire_man_prod_w_lg_w_vector2_range4899w4900w(0) <= wire_man_prod_w_vector2_range4899w(0) XOR wire_man_prod_w_neg_msb_range3779w(0);
	wire_man_prod_w_lg_w_vector2_range4909w4910w(0) <= wire_man_prod_w_vector2_range4909w(0) XOR wire_man_prod_w_neg_msb_range3775w(0);
	wire_man_prod_w_lg_w_vector2_range4919w4920w(0) <= wire_man_prod_w_vector2_range4919w(0) XOR wire_man_prod_w_neg_msb_range3771w(0);
	wire_man_prod_w_lg_w_vector2_range4929w4930w(0) <= wire_man_prod_w_vector2_range4929w(0) XOR wire_man_prod_w_neg_msb_range3767w(0);
	wire_man_prod_w_lg_w_vector2_range4939w4940w(0) <= wire_man_prod_w_vector2_range4939w(0) XOR wire_man_prod_w_neg_msb_range3763w(0);
	wire_man_prod_w_lg_w_vector2_range4949w4950w(0) <= wire_man_prod_w_vector2_range4949w(0) XOR wire_man_prod_w_neg_msb_range3759w(0);
	wire_man_prod_w_lg_w_vector2_range4959w4960w(0) <= wire_man_prod_w_vector2_range4959w(0) XOR wire_man_prod_w_neg_msb_range3755w(0);
	wire_man_prod_w_lg_w_vector2_range4969w4970w(0) <= wire_man_prod_w_vector2_range4969w(0) XOR wire_man_prod_w_neg_msb_range3751w(0);
	wire_man_prod_w_lg_w_vector2_range4979w4980w(0) <= wire_man_prod_w_vector2_range4979w(0) XOR wire_man_prod_w_neg_msb_range3747w(0);
	wire_man_prod_w_lg_w_vector2_range4259w4260w(0) <= wire_man_prod_w_vector2_range4259w(0) XOR wire_man_prod_w_neg_msb_range4141w(0);
	wire_man_prod_w_lg_w_vector2_range4989w4990w(0) <= wire_man_prod_w_vector2_range4989w(0) XOR wire_man_prod_w_neg_msb_range3743w(0);
	wire_man_prod_w_lg_w_vector2_range4999w5000w(0) <= wire_man_prod_w_vector2_range4999w(0) XOR wire_man_prod_w_neg_msb_range3739w(0);
	wire_man_prod_w_lg_w_vector2_range5009w5010w(0) <= wire_man_prod_w_vector2_range5009w(0) XOR wire_man_prod_w_neg_msb_range3735w(0);
	wire_man_prod_w_lg_w_vector2_range5019w5020w(0) <= wire_man_prod_w_vector2_range5019w(0) XOR wire_man_prod_w_neg_msb_range3731w(0);
	wire_man_prod_w_lg_w_vector2_range5029w5030w(0) <= wire_man_prod_w_vector2_range5029w(0) XOR wire_man_prod_w_neg_msb_range3727w(0);
	wire_man_prod_w_lg_w_vector2_range5039w5040w(0) <= wire_man_prod_w_vector2_range5039w(0) XOR wire_man_prod_w_neg_msb_range3723w(0);
	wire_man_prod_w_lg_w_vector2_range5049w5050w(0) <= wire_man_prod_w_vector2_range5049w(0) XOR wire_man_prod_w_neg_msb_range3719w(0);
	wire_man_prod_w_lg_w_vector2_range5059w5060w(0) <= wire_man_prod_w_vector2_range5059w(0) XOR wire_man_prod_w_neg_msb_range3715w(0);
	wire_man_prod_w_lg_w_vector2_range5069w5070w(0) <= wire_man_prod_w_vector2_range5069w(0) XOR wire_man_prod_w_neg_msb_range3711w(0);
	wire_man_prod_w_lg_w_vector2_range5079w5080w(0) <= wire_man_prod_w_vector2_range5079w(0) XOR wire_man_prod_w_neg_msb_range3705w(0);
	wire_man_prod_w_lg_w_vector2_range4269w4270w(0) <= wire_man_prod_w_vector2_range4269w(0) XOR wire_man_prod_w_neg_msb_range4135w(0);
	wire_man_prod_w_lg_w_vector2_range4279w4280w(0) <= wire_man_prod_w_vector2_range4279w(0) XOR wire_man_prod_w_neg_msb_range4129w(0);
	car_one <= ( wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5079w5085w5086w5087w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5069w5075w5076w5077w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5059w5065w5066w5067w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5049w5055w5056w5057w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5039w5045w5046w5047w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5029w5035w5036w5037w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5019w5025w5026w5027w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range5009w5015w5016w5017w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4999w5005w5006w5007w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4989w4995w4996w4997w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4979w4985w4986w4987w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4969w4975w4976w4977w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4959w4965w4966w4967w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4949w4955w4956w4957w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4939w4945w4946w4947w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4929w4935w4936w4937w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4919w4925w4926w4927w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4909w4915w4916w4917w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4899w4905w4906w4907w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4889w4895w4896w4897w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4879w4885w4886w4887w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4869w4875w4876w4877w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4859w4865w4866w4867w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4849w4855w4856w4857w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4839w4845w4846w4847w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4829w4835w4836w4837w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4819w4825w4826w4827w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4809w4815w4816w4817w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4799w4805w4806w4807w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4789w4795w4796w4797w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4779w4785w4786w4787w
 & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4769w4775w4776w4777w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4759w4765w4766w4767w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4749w4755w4756w4757w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4739w4745w4746w4747w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4729w4735w4736w4737w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4719w4725w4726w4727w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4709w4715w4716w4717w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4699w4705w4706w4707w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4689w4695w4696w4697w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4679w4685w4686w4687w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4669w4675w4676w4677w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4659w4665w4666w4667w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4649w4655w4656w4657w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4639w4645w4646w4647w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4629w4635w4636w4637w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4619w4625w4626w4627w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4609w4615w4616w4617w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4599w4605w4606w4607w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4589w4595w4596w4597w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4579w4585w4586w4587w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4569w4575w4576w4577w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4559w4565w4566w4567w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4549w4555w4556w4557w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4539w4545w4546w4547w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4529w4535w4536w4537w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4519w4525w4526w4527w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4509w4515w4516w4517w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4499w4505w4506w4507w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4489w4495w4496w4497w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4479w4485w4486w4487w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4469w4475w4476w4477w
 & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4459w4465w4466w4467w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4449w4455w4456w4457w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4439w4445w4446w4447w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4429w4435w4436w4437w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4419w4425w4426w4427w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4409w4415w4416w4417w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4399w4405w4406w4407w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4389w4395w4396w4397w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4379w4385w4386w4387w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4369w4375w4376w4377w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4359w4365w4366w4367w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4349w4355w4356w4357w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4339w4345w4346w4347w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4329w4335w4336w4337w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4319w4325w4326w4327w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4309w4315w4316w4317w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4299w4305w4306w4307w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4289w4295w4296w4297w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4279w4285w4286w4287w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4269w4275w4276w4277w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4259w4265w4266w4267w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4249w4255w4256w4257w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4239w4245w4246w4247w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4229w4235w4236w4237w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4219w4225w4226w4227w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4209w4215w4216w4217w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4199w4205w4206w4207w & wire_man_prod_w_lg_w_lg_w_lg_w_vector2_range4187w4194w4195w4196w);
	car_one_adj <= ( car_one(88 DOWNTO 0) & "1");
	car_two <= ( wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6075w6081w6082w6083w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6064w6070w6071w6072w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6053w6059w6060w6061w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6042w6048w6049w6050w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6031w6037w6038w6039w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6020w6026w6027w6028w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range6009w6015w6016w6017w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5998w6004w6005w6006w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5987w5993w5994w5995w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5976w5982w5983w5984w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5965w5971w5972w5973w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5954w5960w5961w5962w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5943w5949w5950w5951w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5932w5938w5939w5940w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5921w5927w5928w5929w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5910w5916w5917w5918w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5899w5905w5906w5907w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5888w5894w5895w5896w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5877w5883w5884w5885w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5866w5872w5873w5874w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5855w5861w5862w5863w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5844w5850w5851w5852w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5833w5839w5840w5841w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5822w5828w5829w5830w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5811w5817w5818w5819w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5800w5806w5807w5808w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5789w5795w5796w5797w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5778w5784w5785w5786w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5767w5773w5774w5775w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5756w5762w5763w5764w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5745w5751w5752w5753w
 & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5734w5740w5741w5742w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5723w5729w5730w5731w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5712w5718w5719w5720w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5701w5707w5708w5709w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5690w5696w5697w5698w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5679w5685w5686w5687w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5668w5674w5675w5676w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5657w5663w5664w5665w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5646w5652w5653w5654w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5635w5641w5642w5643w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5624w5630w5631w5632w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5613w5619w5620w5621w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5602w5608w5609w5610w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5591w5597w5598w5599w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5580w5586w5587w5588w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5569w5575w5576w5577w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5558w5564w5565w5566w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5547w5553w5554w5555w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5536w5542w5543w5544w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5525w5531w5532w5533w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5514w5520w5521w5522w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5503w5509w5510w5511w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5492w5498w5499w5500w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5481w5487w5488w5489w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5470w5476w5477w5478w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5459w5465w5466w5467w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5448w5454w5455w5456w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5437w5443w5444w5445w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5426w5432w5433w5434w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5415w5421w5422w5423w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5404w5410w5411w5412w
 & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5393w5399w5400w5401w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5382w5388w5389w5390w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5371w5377w5378w5379w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5360w5366w5367w5368w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5349w5355w5356w5357w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5338w5344w5345w5346w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5327w5333w5334w5335w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5316w5322w5323w5324w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5305w5311w5312w5313w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5294w5300w5301w5302w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5283w5289w5290w5291w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5272w5278w5279w5280w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5261w5267w5268w5269w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5250w5256w5257w5258w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5239w5245w5246w5247w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5228w5234w5235w5236w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5217w5223w5224w5225w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5206w5212w5213w5214w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5195w5201w5202w5203w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5184w5190w5191w5192w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5173w5179w5180w5181w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5162w5168w5169w5170w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5151w5157w5158w5159w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5140w5146w5147w5148w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5129w5135w5136w5137w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5118w5124w5125w5126w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5107w5113w5114w5115w & wire_man_prod_w_lg_w_lg_w_lg_w_vector1_range5094w5101w5102w5103w);
	car_two_adj <= ( car_two(88 DOWNTO 0) & "1");
	car_two_wo <= car_two_adj_reg0;
	lowest_bits_wi <= lsb_prod_wo(29 DOWNTO 0);
	lowest_bits_wo <= lowest_bits_wi_reg1;
	lsb_prod_wi <= wire_lsb_prod_result;
	lsb_prod_wo <= lsb_prod_wi_reg0;
	mid_prod_wi <= wire_mid_prod_result;
	mid_prod_wo <= mid_prod_wi_reg0;
	msb_prod_out <= wire_msb_prod_result;
	msb_prod_wi <= msb_prod_out;
	msb_prod_wo <= msb_prod_wi_reg0;
	neg_lsb <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & wire_man_prod_w_lg_w_lsb_prod_wo_range3830w3831w & wire_man_prod_w_lg_w_lsb_prod_wo_range3836w3837w & wire_man_prod_w_lg_w_lsb_prod_wo_range3842w3843w & wire_man_prod_w_lg_w_lsb_prod_wo_range3848w3849w & wire_man_prod_w_lg_w_lsb_prod_wo_range3854w3855w & wire_man_prod_w_lg_w_lsb_prod_wo_range3860w3861w & wire_man_prod_w_lg_w_lsb_prod_wo_range3866w3867w & wire_man_prod_w_lg_w_lsb_prod_wo_range3872w3873w & wire_man_prod_w_lg_w_lsb_prod_wo_range3878w3879w & wire_man_prod_w_lg_w_lsb_prod_wo_range3884w3885w & wire_man_prod_w_lg_w_lsb_prod_wo_range3890w3891w & wire_man_prod_w_lg_w_lsb_prod_wo_range3896w3897w & wire_man_prod_w_lg_w_lsb_prod_wo_range3902w3903w & wire_man_prod_w_lg_w_lsb_prod_wo_range3908w3909w & wire_man_prod_w_lg_w_lsb_prod_wo_range3914w3915w & wire_man_prod_w_lg_w_lsb_prod_wo_range3920w3921w & wire_man_prod_w_lg_w_lsb_prod_wo_range3926w3927w & wire_man_prod_w_lg_w_lsb_prod_wo_range3932w3933w & wire_man_prod_w_lg_w_lsb_prod_wo_range3938w3939w & wire_man_prod_w_lg_w_lsb_prod_wo_range3944w3945w & wire_man_prod_w_lg_w_lsb_prod_wo_range3950w3951w & wire_man_prod_w_lg_w_lsb_prod_wo_range3956w3957w & wire_man_prod_w_lg_w_lsb_prod_wo_range3962w3963w & wire_man_prod_w_lg_w_lsb_prod_wo_range3968w3969w & wire_man_prod_w_lg_w_lsb_prod_wo_range3974w3975w & wire_man_prod_w_lg_w_lsb_prod_wo_range3980w3981w & wire_man_prod_w_lg_w_lsb_prod_wo_range3986w3987w & wire_man_prod_w_lg_w_lsb_prod_wo_range3992w3993w & wire_man_prod_w_lg_w_lsb_prod_wo_range3998w3999w & wire_man_prod_w_lg_w_lsb_prod_wo_range4004w4005w & wire_man_prod_w_lg_w_lsb_prod_wo_range4010w4011w & wire_man_prod_w_lg_w_lsb_prod_wo_range4016w4017w & wire_man_prod_w_lg_w_lsb_prod_wo_range4022w4023w & wire_man_prod_w_lg_w_lsb_prod_wo_range4028w4029w & wire_man_prod_w_lg_w_lsb_prod_wo_range4034w4035w & wire_man_prod_w_lg_w_lsb_prod_wo_range4040w4041w & wire_man_prod_w_lg_w_lsb_prod_wo_range4046w4047w
 & wire_man_prod_w_lg_w_lsb_prod_wo_range4052w4053w & wire_man_prod_w_lg_w_lsb_prod_wo_range4058w4059w & wire_man_prod_w_lg_w_lsb_prod_wo_range4064w4065w & wire_man_prod_w_lg_w_lsb_prod_wo_range4070w4071w & wire_man_prod_w_lg_w_lsb_prod_wo_range4076w4077w & wire_man_prod_w_lg_w_lsb_prod_wo_range4082w4083w & wire_man_prod_w_lg_w_lsb_prod_wo_range4088w4089w & wire_man_prod_w_lg_w_lsb_prod_wo_range4094w4095w & wire_man_prod_w_lg_w_lsb_prod_wo_range4100w4101w & wire_man_prod_w_lg_w_lsb_prod_wo_range4106w4107w & wire_man_prod_w_lg_w_lsb_prod_wo_range4112w4113w & wire_man_prod_w_lg_w_lsb_prod_wo_range4118w4119w & wire_man_prod_w_lg_w_lsb_prod_wo_range4124w4125w & wire_man_prod_w_lg_w_lsb_prod_wo_range4130w4131w & wire_man_prod_w_lg_w_lsb_prod_wo_range4136w4137w & wire_man_prod_w_lg_w_lsb_prod_wo_range4142w4143w & wire_man_prod_w_lg_w_lsb_prod_wo_range4148w4149w & wire_man_prod_w_lg_w_lsb_prod_wo_range4154w4155w & wire_man_prod_w_lg_w_lsb_prod_wo_range4160w4161w & wire_man_prod_w_lg_w_lsb_prod_wo_range4166w4167w & wire_man_prod_w_lg_w_lsb_prod_wo_range4172w4173w & wire_man_prod_w_lg_w_lsb_prod_wo_range4178w4179w & wire_man_prod_w_lg_w_lsb_prod_wo_range4184w4185w);
	neg_msb <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & wire_man_prod_w_lg_w_msb_prod_wo_range3827w3828w & wire_man_prod_w_lg_w_msb_prod_wo_range3833w3834w & wire_man_prod_w_lg_w_msb_prod_wo_range3839w3840w & wire_man_prod_w_lg_w_msb_prod_wo_range3845w3846w & wire_man_prod_w_lg_w_msb_prod_wo_range3851w3852w & wire_man_prod_w_lg_w_msb_prod_wo_range3857w3858w & wire_man_prod_w_lg_w_msb_prod_wo_range3863w3864w & wire_man_prod_w_lg_w_msb_prod_wo_range3869w3870w & wire_man_prod_w_lg_w_msb_prod_wo_range3875w3876w & wire_man_prod_w_lg_w_msb_prod_wo_range3881w3882w & wire_man_prod_w_lg_w_msb_prod_wo_range3887w3888w & wire_man_prod_w_lg_w_msb_prod_wo_range3893w3894w & wire_man_prod_w_lg_w_msb_prod_wo_range3899w3900w & wire_man_prod_w_lg_w_msb_prod_wo_range3905w3906w & wire_man_prod_w_lg_w_msb_prod_wo_range3911w3912w & wire_man_prod_w_lg_w_msb_prod_wo_range3917w3918w & wire_man_prod_w_lg_w_msb_prod_wo_range3923w3924w & wire_man_prod_w_lg_w_msb_prod_wo_range3929w3930w & wire_man_prod_w_lg_w_msb_prod_wo_range3935w3936w & wire_man_prod_w_lg_w_msb_prod_wo_range3941w3942w & wire_man_prod_w_lg_w_msb_prod_wo_range3947w3948w & wire_man_prod_w_lg_w_msb_prod_wo_range3953w3954w & wire_man_prod_w_lg_w_msb_prod_wo_range3959w3960w & wire_man_prod_w_lg_w_msb_prod_wo_range3965w3966w & wire_man_prod_w_lg_w_msb_prod_wo_range3971w3972w & wire_man_prod_w_lg_w_msb_prod_wo_range3977w3978w & wire_man_prod_w_lg_w_msb_prod_wo_range3983w3984w & wire_man_prod_w_lg_w_msb_prod_wo_range3989w3990w & wire_man_prod_w_lg_w_msb_prod_wo_range3995w3996w & wire_man_prod_w_lg_w_msb_prod_wo_range4001w4002w & wire_man_prod_w_lg_w_msb_prod_wo_range4007w4008w & wire_man_prod_w_lg_w_msb_prod_wo_range4013w4014w & wire_man_prod_w_lg_w_msb_prod_wo_range4019w4020w & wire_man_prod_w_lg_w_msb_prod_wo_range4025w4026w & wire_man_prod_w_lg_w_msb_prod_wo_range4031w4032w & wire_man_prod_w_lg_w_msb_prod_wo_range4037w4038w & wire_man_prod_w_lg_w_msb_prod_wo_range4043w4044w
 & wire_man_prod_w_lg_w_msb_prod_wo_range4049w4050w & wire_man_prod_w_lg_w_msb_prod_wo_range4055w4056w & wire_man_prod_w_lg_w_msb_prod_wo_range4061w4062w & wire_man_prod_w_lg_w_msb_prod_wo_range4067w4068w & wire_man_prod_w_lg_w_msb_prod_wo_range4073w4074w & wire_man_prod_w_lg_w_msb_prod_wo_range4079w4080w & wire_man_prod_w_lg_w_msb_prod_wo_range4085w4086w & wire_man_prod_w_lg_w_msb_prod_wo_range4091w4092w & wire_man_prod_w_lg_w_msb_prod_wo_range4097w4098w & wire_man_prod_w_lg_w_msb_prod_wo_range4103w4104w & wire_man_prod_w_lg_w_msb_prod_wo_range4109w4110w & wire_man_prod_w_lg_w_msb_prod_wo_range4115w4116w & wire_man_prod_w_lg_w_msb_prod_wo_range4121w4122w & wire_man_prod_w_lg_w_msb_prod_wo_range4127w4128w & wire_man_prod_w_lg_w_msb_prod_wo_range4133w4134w & wire_man_prod_w_lg_w_msb_prod_wo_range4139w4140w & wire_man_prod_w_lg_w_msb_prod_wo_range4145w4146w & wire_man_prod_w_lg_w_msb_prod_wo_range4151w4152w & wire_man_prod_w_lg_w_msb_prod_wo_range4157w4158w & wire_man_prod_w_lg_w_msb_prod_wo_range4163w4164w & wire_man_prod_w_lg_w_msb_prod_wo_range4169w4170w & wire_man_prod_w_lg_w_msb_prod_wo_range4175w4176w & wire_man_prod_w_lg_w_msb_prod_wo_range4181w4182w);
	result <= ( wire_sum_result(89 DOWNTO 0) & lowest_bits_wo);
	sum_one <= ( wire_man_prod_w_lg_w_lg_w_vector2_range5079w5080w5081w & wire_man_prod_w_lg_w_lg_w_vector2_range5069w5070w5071w & wire_man_prod_w_lg_w_lg_w_vector2_range5059w5060w5061w & wire_man_prod_w_lg_w_lg_w_vector2_range5049w5050w5051w & wire_man_prod_w_lg_w_lg_w_vector2_range5039w5040w5041w & wire_man_prod_w_lg_w_lg_w_vector2_range5029w5030w5031w & wire_man_prod_w_lg_w_lg_w_vector2_range5019w5020w5021w & wire_man_prod_w_lg_w_lg_w_vector2_range5009w5010w5011w & wire_man_prod_w_lg_w_lg_w_vector2_range4999w5000w5001w & wire_man_prod_w_lg_w_lg_w_vector2_range4989w4990w4991w & wire_man_prod_w_lg_w_lg_w_vector2_range4979w4980w4981w & wire_man_prod_w_lg_w_lg_w_vector2_range4969w4970w4971w & wire_man_prod_w_lg_w_lg_w_vector2_range4959w4960w4961w & wire_man_prod_w_lg_w_lg_w_vector2_range4949w4950w4951w & wire_man_prod_w_lg_w_lg_w_vector2_range4939w4940w4941w & wire_man_prod_w_lg_w_lg_w_vector2_range4929w4930w4931w & wire_man_prod_w_lg_w_lg_w_vector2_range4919w4920w4921w & wire_man_prod_w_lg_w_lg_w_vector2_range4909w4910w4911w & wire_man_prod_w_lg_w_lg_w_vector2_range4899w4900w4901w & wire_man_prod_w_lg_w_lg_w_vector2_range4889w4890w4891w & wire_man_prod_w_lg_w_lg_w_vector2_range4879w4880w4881w & wire_man_prod_w_lg_w_lg_w_vector2_range4869w4870w4871w & wire_man_prod_w_lg_w_lg_w_vector2_range4859w4860w4861w & wire_man_prod_w_lg_w_lg_w_vector2_range4849w4850w4851w & wire_man_prod_w_lg_w_lg_w_vector2_range4839w4840w4841w & wire_man_prod_w_lg_w_lg_w_vector2_range4829w4830w4831w & wire_man_prod_w_lg_w_lg_w_vector2_range4819w4820w4821w & wire_man_prod_w_lg_w_lg_w_vector2_range4809w4810w4811w & wire_man_prod_w_lg_w_lg_w_vector2_range4799w4800w4801w & wire_man_prod_w_lg_w_lg_w_vector2_range4789w4790w4791w & wire_man_prod_w_lg_w_lg_w_vector2_range4779w4780w4781w & wire_man_prod_w_lg_w_lg_w_vector2_range4769w4770w4771w & wire_man_prod_w_lg_w_lg_w_vector2_range4759w4760w4761w & wire_man_prod_w_lg_w_lg_w_vector2_range4749w4750w4751w & wire_man_prod_w_lg_w_lg_w_vector2_range4739w4740w4741w & wire_man_prod_w_lg_w_lg_w_vector2_range4729w4730w4731w
 & wire_man_prod_w_lg_w_lg_w_vector2_range4719w4720w4721w & wire_man_prod_w_lg_w_lg_w_vector2_range4709w4710w4711w & wire_man_prod_w_lg_w_lg_w_vector2_range4699w4700w4701w & wire_man_prod_w_lg_w_lg_w_vector2_range4689w4690w4691w & wire_man_prod_w_lg_w_lg_w_vector2_range4679w4680w4681w & wire_man_prod_w_lg_w_lg_w_vector2_range4669w4670w4671w & wire_man_prod_w_lg_w_lg_w_vector2_range4659w4660w4661w & wire_man_prod_w_lg_w_lg_w_vector2_range4649w4650w4651w & wire_man_prod_w_lg_w_lg_w_vector2_range4639w4640w4641w & wire_man_prod_w_lg_w_lg_w_vector2_range4629w4630w4631w & wire_man_prod_w_lg_w_lg_w_vector2_range4619w4620w4621w & wire_man_prod_w_lg_w_lg_w_vector2_range4609w4610w4611w & wire_man_prod_w_lg_w_lg_w_vector2_range4599w4600w4601w & wire_man_prod_w_lg_w_lg_w_vector2_range4589w4590w4591w & wire_man_prod_w_lg_w_lg_w_vector2_range4579w4580w4581w & wire_man_prod_w_lg_w_lg_w_vector2_range4569w4570w4571w & wire_man_prod_w_lg_w_lg_w_vector2_range4559w4560w4561w & wire_man_prod_w_lg_w_lg_w_vector2_range4549w4550w4551w & wire_man_prod_w_lg_w_lg_w_vector2_range4539w4540w4541w & wire_man_prod_w_lg_w_lg_w_vector2_range4529w4530w4531w & wire_man_prod_w_lg_w_lg_w_vector2_range4519w4520w4521w & wire_man_prod_w_lg_w_lg_w_vector2_range4509w4510w4511w & wire_man_prod_w_lg_w_lg_w_vector2_range4499w4500w4501w & wire_man_prod_w_lg_w_lg_w_vector2_range4489w4490w4491w & wire_man_prod_w_lg_w_lg_w_vector2_range4479w4480w4481w & wire_man_prod_w_lg_w_lg_w_vector2_range4469w4470w4471w & wire_man_prod_w_lg_w_lg_w_vector2_range4459w4460w4461w & wire_man_prod_w_lg_w_lg_w_vector2_range4449w4450w4451w & wire_man_prod_w_lg_w_lg_w_vector2_range4439w4440w4441w & wire_man_prod_w_lg_w_lg_w_vector2_range4429w4430w4431w & wire_man_prod_w_lg_w_lg_w_vector2_range4419w4420w4421w & wire_man_prod_w_lg_w_lg_w_vector2_range4409w4410w4411w & wire_man_prod_w_lg_w_lg_w_vector2_range4399w4400w4401w & wire_man_prod_w_lg_w_lg_w_vector2_range4389w4390w4391w & wire_man_prod_w_lg_w_lg_w_vector2_range4379w4380w4381w & wire_man_prod_w_lg_w_lg_w_vector2_range4369w4370w4371w
 & wire_man_prod_w_lg_w_lg_w_vector2_range4359w4360w4361w & wire_man_prod_w_lg_w_lg_w_vector2_range4349w4350w4351w & wire_man_prod_w_lg_w_lg_w_vector2_range4339w4340w4341w & wire_man_prod_w_lg_w_lg_w_vector2_range4329w4330w4331w & wire_man_prod_w_lg_w_lg_w_vector2_range4319w4320w4321w & wire_man_prod_w_lg_w_lg_w_vector2_range4309w4310w4311w & wire_man_prod_w_lg_w_lg_w_vector2_range4299w4300w4301w & wire_man_prod_w_lg_w_lg_w_vector2_range4289w4290w4291w & wire_man_prod_w_lg_w_lg_w_vector2_range4279w4280w4281w & wire_man_prod_w_lg_w_lg_w_vector2_range4269w4270w4271w & wire_man_prod_w_lg_w_lg_w_vector2_range4259w4260w4261w & wire_man_prod_w_lg_w_lg_w_vector2_range4249w4250w4251w & wire_man_prod_w_lg_w_lg_w_vector2_range4239w4240w4241w & wire_man_prod_w_lg_w_lg_w_vector2_range4229w4230w4231w & wire_man_prod_w_lg_w_lg_w_vector2_range4219w4220w4221w & wire_man_prod_w_lg_w_lg_w_vector2_range4209w4210w4211w & wire_man_prod_w_lg_w_lg_w_vector2_range4199w4200w4201w & wire_man_prod_w_lg_w_lg_w_vector2_range4187w4188w4189w);
	sum_two <= ( wire_man_prod_w_lg_w_lg_w_vector1_range6075w6076w6077w & wire_man_prod_w_lg_w_lg_w_vector1_range6064w6065w6066w & wire_man_prod_w_lg_w_lg_w_vector1_range6053w6054w6055w & wire_man_prod_w_lg_w_lg_w_vector1_range6042w6043w6044w & wire_man_prod_w_lg_w_lg_w_vector1_range6031w6032w6033w & wire_man_prod_w_lg_w_lg_w_vector1_range6020w6021w6022w & wire_man_prod_w_lg_w_lg_w_vector1_range6009w6010w6011w & wire_man_prod_w_lg_w_lg_w_vector1_range5998w5999w6000w & wire_man_prod_w_lg_w_lg_w_vector1_range5987w5988w5989w & wire_man_prod_w_lg_w_lg_w_vector1_range5976w5977w5978w & wire_man_prod_w_lg_w_lg_w_vector1_range5965w5966w5967w & wire_man_prod_w_lg_w_lg_w_vector1_range5954w5955w5956w & wire_man_prod_w_lg_w_lg_w_vector1_range5943w5944w5945w & wire_man_prod_w_lg_w_lg_w_vector1_range5932w5933w5934w & wire_man_prod_w_lg_w_lg_w_vector1_range5921w5922w5923w & wire_man_prod_w_lg_w_lg_w_vector1_range5910w5911w5912w & wire_man_prod_w_lg_w_lg_w_vector1_range5899w5900w5901w & wire_man_prod_w_lg_w_lg_w_vector1_range5888w5889w5890w & wire_man_prod_w_lg_w_lg_w_vector1_range5877w5878w5879w & wire_man_prod_w_lg_w_lg_w_vector1_range5866w5867w5868w & wire_man_prod_w_lg_w_lg_w_vector1_range5855w5856w5857w & wire_man_prod_w_lg_w_lg_w_vector1_range5844w5845w5846w & wire_man_prod_w_lg_w_lg_w_vector1_range5833w5834w5835w & wire_man_prod_w_lg_w_lg_w_vector1_range5822w5823w5824w & wire_man_prod_w_lg_w_lg_w_vector1_range5811w5812w5813w & wire_man_prod_w_lg_w_lg_w_vector1_range5800w5801w5802w & wire_man_prod_w_lg_w_lg_w_vector1_range5789w5790w5791w & wire_man_prod_w_lg_w_lg_w_vector1_range5778w5779w5780w & wire_man_prod_w_lg_w_lg_w_vector1_range5767w5768w5769w & wire_man_prod_w_lg_w_lg_w_vector1_range5756w5757w5758w & wire_man_prod_w_lg_w_lg_w_vector1_range5745w5746w5747w & wire_man_prod_w_lg_w_lg_w_vector1_range5734w5735w5736w & wire_man_prod_w_lg_w_lg_w_vector1_range5723w5724w5725w & wire_man_prod_w_lg_w_lg_w_vector1_range5712w5713w5714w & wire_man_prod_w_lg_w_lg_w_vector1_range5701w5702w5703w & wire_man_prod_w_lg_w_lg_w_vector1_range5690w5691w5692w
 & wire_man_prod_w_lg_w_lg_w_vector1_range5679w5680w5681w & wire_man_prod_w_lg_w_lg_w_vector1_range5668w5669w5670w & wire_man_prod_w_lg_w_lg_w_vector1_range5657w5658w5659w & wire_man_prod_w_lg_w_lg_w_vector1_range5646w5647w5648w & wire_man_prod_w_lg_w_lg_w_vector1_range5635w5636w5637w & wire_man_prod_w_lg_w_lg_w_vector1_range5624w5625w5626w & wire_man_prod_w_lg_w_lg_w_vector1_range5613w5614w5615w & wire_man_prod_w_lg_w_lg_w_vector1_range5602w5603w5604w & wire_man_prod_w_lg_w_lg_w_vector1_range5591w5592w5593w & wire_man_prod_w_lg_w_lg_w_vector1_range5580w5581w5582w & wire_man_prod_w_lg_w_lg_w_vector1_range5569w5570w5571w & wire_man_prod_w_lg_w_lg_w_vector1_range5558w5559w5560w & wire_man_prod_w_lg_w_lg_w_vector1_range5547w5548w5549w & wire_man_prod_w_lg_w_lg_w_vector1_range5536w5537w5538w & wire_man_prod_w_lg_w_lg_w_vector1_range5525w5526w5527w & wire_man_prod_w_lg_w_lg_w_vector1_range5514w5515w5516w & wire_man_prod_w_lg_w_lg_w_vector1_range5503w5504w5505w & wire_man_prod_w_lg_w_lg_w_vector1_range5492w5493w5494w & wire_man_prod_w_lg_w_lg_w_vector1_range5481w5482w5483w & wire_man_prod_w_lg_w_lg_w_vector1_range5470w5471w5472w & wire_man_prod_w_lg_w_lg_w_vector1_range5459w5460w5461w & wire_man_prod_w_lg_w_lg_w_vector1_range5448w5449w5450w & wire_man_prod_w_lg_w_lg_w_vector1_range5437w5438w5439w & wire_man_prod_w_lg_w_lg_w_vector1_range5426w5427w5428w & wire_man_prod_w_lg_w_lg_w_vector1_range5415w5416w5417w & wire_man_prod_w_lg_w_lg_w_vector1_range5404w5405w5406w & wire_man_prod_w_lg_w_lg_w_vector1_range5393w5394w5395w & wire_man_prod_w_lg_w_lg_w_vector1_range5382w5383w5384w & wire_man_prod_w_lg_w_lg_w_vector1_range5371w5372w5373w & wire_man_prod_w_lg_w_lg_w_vector1_range5360w5361w5362w & wire_man_prod_w_lg_w_lg_w_vector1_range5349w5350w5351w & wire_man_prod_w_lg_w_lg_w_vector1_range5338w5339w5340w & wire_man_prod_w_lg_w_lg_w_vector1_range5327w5328w5329w & wire_man_prod_w_lg_w_lg_w_vector1_range5316w5317w5318w & wire_man_prod_w_lg_w_lg_w_vector1_range5305w5306w5307w & wire_man_prod_w_lg_w_lg_w_vector1_range5294w5295w5296w
 & wire_man_prod_w_lg_w_lg_w_vector1_range5283w5284w5285w & wire_man_prod_w_lg_w_lg_w_vector1_range5272w5273w5274w & wire_man_prod_w_lg_w_lg_w_vector1_range5261w5262w5263w & wire_man_prod_w_lg_w_lg_w_vector1_range5250w5251w5252w & wire_man_prod_w_lg_w_lg_w_vector1_range5239w5240w5241w & wire_man_prod_w_lg_w_lg_w_vector1_range5228w5229w5230w & wire_man_prod_w_lg_w_lg_w_vector1_range5217w5218w5219w & wire_man_prod_w_lg_w_lg_w_vector1_range5206w5207w5208w & wire_man_prod_w_lg_w_lg_w_vector1_range5195w5196w5197w & wire_man_prod_w_lg_w_lg_w_vector1_range5184w5185w5186w & wire_man_prod_w_lg_w_lg_w_vector1_range5173w5174w5175w & wire_man_prod_w_lg_w_lg_w_vector1_range5162w5163w5164w & wire_man_prod_w_lg_w_lg_w_vector1_range5151w5152w5153w & wire_man_prod_w_lg_w_lg_w_vector1_range5140w5141w5142w & wire_man_prod_w_lg_w_lg_w_vector1_range5129w5130w5131w & wire_man_prod_w_lg_w_lg_w_vector1_range5118w5119w5120w & wire_man_prod_w_lg_w_lg_w_vector1_range5107w5108w5109w & wire_man_prod_w_lg_w_lg_w_vector1_range5094w5095w5096w);
	sum_two_wo <= sum_two_reg0;
	vector1 <= ( msb_prod_wo & lsb_prod_wo(59 DOWNTO 30));
	vector2 <= ( "0000000000000000000000000000" & mid_prod_wo);
	wire_a <= dataa;
	wire_b <= datab;
	wire_man_prod_w_car_one_adj_range5092w(0) <= car_one_adj(0);
	wire_man_prod_w_car_one_adj_range5205w(0) <= car_one_adj(10);
	wire_man_prod_w_car_one_adj_range5216w(0) <= car_one_adj(11);
	wire_man_prod_w_car_one_adj_range5227w(0) <= car_one_adj(12);
	wire_man_prod_w_car_one_adj_range5238w(0) <= car_one_adj(13);
	wire_man_prod_w_car_one_adj_range5249w(0) <= car_one_adj(14);
	wire_man_prod_w_car_one_adj_range5260w(0) <= car_one_adj(15);
	wire_man_prod_w_car_one_adj_range5271w(0) <= car_one_adj(16);
	wire_man_prod_w_car_one_adj_range5282w(0) <= car_one_adj(17);
	wire_man_prod_w_car_one_adj_range5293w(0) <= car_one_adj(18);
	wire_man_prod_w_car_one_adj_range5304w(0) <= car_one_adj(19);
	wire_man_prod_w_car_one_adj_range5106w(0) <= car_one_adj(1);
	wire_man_prod_w_car_one_adj_range5315w(0) <= car_one_adj(20);
	wire_man_prod_w_car_one_adj_range5326w(0) <= car_one_adj(21);
	wire_man_prod_w_car_one_adj_range5337w(0) <= car_one_adj(22);
	wire_man_prod_w_car_one_adj_range5348w(0) <= car_one_adj(23);
	wire_man_prod_w_car_one_adj_range5359w(0) <= car_one_adj(24);
	wire_man_prod_w_car_one_adj_range5370w(0) <= car_one_adj(25);
	wire_man_prod_w_car_one_adj_range5381w(0) <= car_one_adj(26);
	wire_man_prod_w_car_one_adj_range5392w(0) <= car_one_adj(27);
	wire_man_prod_w_car_one_adj_range5403w(0) <= car_one_adj(28);
	wire_man_prod_w_car_one_adj_range5414w(0) <= car_one_adj(29);
	wire_man_prod_w_car_one_adj_range5117w(0) <= car_one_adj(2);
	wire_man_prod_w_car_one_adj_range5425w(0) <= car_one_adj(30);
	wire_man_prod_w_car_one_adj_range5436w(0) <= car_one_adj(31);
	wire_man_prod_w_car_one_adj_range5447w(0) <= car_one_adj(32);
	wire_man_prod_w_car_one_adj_range5458w(0) <= car_one_adj(33);
	wire_man_prod_w_car_one_adj_range5469w(0) <= car_one_adj(34);
	wire_man_prod_w_car_one_adj_range5480w(0) <= car_one_adj(35);
	wire_man_prod_w_car_one_adj_range5491w(0) <= car_one_adj(36);
	wire_man_prod_w_car_one_adj_range5502w(0) <= car_one_adj(37);
	wire_man_prod_w_car_one_adj_range5513w(0) <= car_one_adj(38);
	wire_man_prod_w_car_one_adj_range5524w(0) <= car_one_adj(39);
	wire_man_prod_w_car_one_adj_range5128w(0) <= car_one_adj(3);
	wire_man_prod_w_car_one_adj_range5535w(0) <= car_one_adj(40);
	wire_man_prod_w_car_one_adj_range5546w(0) <= car_one_adj(41);
	wire_man_prod_w_car_one_adj_range5557w(0) <= car_one_adj(42);
	wire_man_prod_w_car_one_adj_range5568w(0) <= car_one_adj(43);
	wire_man_prod_w_car_one_adj_range5579w(0) <= car_one_adj(44);
	wire_man_prod_w_car_one_adj_range5590w(0) <= car_one_adj(45);
	wire_man_prod_w_car_one_adj_range5601w(0) <= car_one_adj(46);
	wire_man_prod_w_car_one_adj_range5612w(0) <= car_one_adj(47);
	wire_man_prod_w_car_one_adj_range5623w(0) <= car_one_adj(48);
	wire_man_prod_w_car_one_adj_range5634w(0) <= car_one_adj(49);
	wire_man_prod_w_car_one_adj_range5139w(0) <= car_one_adj(4);
	wire_man_prod_w_car_one_adj_range5645w(0) <= car_one_adj(50);
	wire_man_prod_w_car_one_adj_range5656w(0) <= car_one_adj(51);
	wire_man_prod_w_car_one_adj_range5667w(0) <= car_one_adj(52);
	wire_man_prod_w_car_one_adj_range5678w(0) <= car_one_adj(53);
	wire_man_prod_w_car_one_adj_range5689w(0) <= car_one_adj(54);
	wire_man_prod_w_car_one_adj_range5700w(0) <= car_one_adj(55);
	wire_man_prod_w_car_one_adj_range5711w(0) <= car_one_adj(56);
	wire_man_prod_w_car_one_adj_range5722w(0) <= car_one_adj(57);
	wire_man_prod_w_car_one_adj_range5733w(0) <= car_one_adj(58);
	wire_man_prod_w_car_one_adj_range5744w(0) <= car_one_adj(59);
	wire_man_prod_w_car_one_adj_range5150w(0) <= car_one_adj(5);
	wire_man_prod_w_car_one_adj_range5755w(0) <= car_one_adj(60);
	wire_man_prod_w_car_one_adj_range5766w(0) <= car_one_adj(61);
	wire_man_prod_w_car_one_adj_range5777w(0) <= car_one_adj(62);
	wire_man_prod_w_car_one_adj_range5788w(0) <= car_one_adj(63);
	wire_man_prod_w_car_one_adj_range5799w(0) <= car_one_adj(64);
	wire_man_prod_w_car_one_adj_range5810w(0) <= car_one_adj(65);
	wire_man_prod_w_car_one_adj_range5821w(0) <= car_one_adj(66);
	wire_man_prod_w_car_one_adj_range5832w(0) <= car_one_adj(67);
	wire_man_prod_w_car_one_adj_range5843w(0) <= car_one_adj(68);
	wire_man_prod_w_car_one_adj_range5854w(0) <= car_one_adj(69);
	wire_man_prod_w_car_one_adj_range5161w(0) <= car_one_adj(6);
	wire_man_prod_w_car_one_adj_range5865w(0) <= car_one_adj(70);
	wire_man_prod_w_car_one_adj_range5876w(0) <= car_one_adj(71);
	wire_man_prod_w_car_one_adj_range5887w(0) <= car_one_adj(72);
	wire_man_prod_w_car_one_adj_range5898w(0) <= car_one_adj(73);
	wire_man_prod_w_car_one_adj_range5909w(0) <= car_one_adj(74);
	wire_man_prod_w_car_one_adj_range5920w(0) <= car_one_adj(75);
	wire_man_prod_w_car_one_adj_range5931w(0) <= car_one_adj(76);
	wire_man_prod_w_car_one_adj_range5942w(0) <= car_one_adj(77);
	wire_man_prod_w_car_one_adj_range5953w(0) <= car_one_adj(78);
	wire_man_prod_w_car_one_adj_range5964w(0) <= car_one_adj(79);
	wire_man_prod_w_car_one_adj_range5172w(0) <= car_one_adj(7);
	wire_man_prod_w_car_one_adj_range5975w(0) <= car_one_adj(80);
	wire_man_prod_w_car_one_adj_range5986w(0) <= car_one_adj(81);
	wire_man_prod_w_car_one_adj_range5997w(0) <= car_one_adj(82);
	wire_man_prod_w_car_one_adj_range6008w(0) <= car_one_adj(83);
	wire_man_prod_w_car_one_adj_range6019w(0) <= car_one_adj(84);
	wire_man_prod_w_car_one_adj_range6030w(0) <= car_one_adj(85);
	wire_man_prod_w_car_one_adj_range6041w(0) <= car_one_adj(86);
	wire_man_prod_w_car_one_adj_range6052w(0) <= car_one_adj(87);
	wire_man_prod_w_car_one_adj_range6063w(0) <= car_one_adj(88);
	wire_man_prod_w_car_one_adj_range6074w(0) <= car_one_adj(89);
	wire_man_prod_w_car_one_adj_range5183w(0) <= car_one_adj(8);
	wire_man_prod_w_car_one_adj_range5194w(0) <= car_one_adj(9);
	wire_man_prod_w_lsb_prod_wo_range4184w(0) <= lsb_prod_wo(0);
	wire_man_prod_w_lsb_prod_wo_range4124w(0) <= lsb_prod_wo(10);
	wire_man_prod_w_lsb_prod_wo_range4118w(0) <= lsb_prod_wo(11);
	wire_man_prod_w_lsb_prod_wo_range4112w(0) <= lsb_prod_wo(12);
	wire_man_prod_w_lsb_prod_wo_range4106w(0) <= lsb_prod_wo(13);
	wire_man_prod_w_lsb_prod_wo_range4100w(0) <= lsb_prod_wo(14);
	wire_man_prod_w_lsb_prod_wo_range4094w(0) <= lsb_prod_wo(15);
	wire_man_prod_w_lsb_prod_wo_range4088w(0) <= lsb_prod_wo(16);
	wire_man_prod_w_lsb_prod_wo_range4082w(0) <= lsb_prod_wo(17);
	wire_man_prod_w_lsb_prod_wo_range4076w(0) <= lsb_prod_wo(18);
	wire_man_prod_w_lsb_prod_wo_range4070w(0) <= lsb_prod_wo(19);
	wire_man_prod_w_lsb_prod_wo_range4178w(0) <= lsb_prod_wo(1);
	wire_man_prod_w_lsb_prod_wo_range4064w(0) <= lsb_prod_wo(20);
	wire_man_prod_w_lsb_prod_wo_range4058w(0) <= lsb_prod_wo(21);
	wire_man_prod_w_lsb_prod_wo_range4052w(0) <= lsb_prod_wo(22);
	wire_man_prod_w_lsb_prod_wo_range4046w(0) <= lsb_prod_wo(23);
	wire_man_prod_w_lsb_prod_wo_range4040w(0) <= lsb_prod_wo(24);
	wire_man_prod_w_lsb_prod_wo_range4034w(0) <= lsb_prod_wo(25);
	wire_man_prod_w_lsb_prod_wo_range4028w(0) <= lsb_prod_wo(26);
	wire_man_prod_w_lsb_prod_wo_range4022w(0) <= lsb_prod_wo(27);
	wire_man_prod_w_lsb_prod_wo_range4016w(0) <= lsb_prod_wo(28);
	wire_man_prod_w_lsb_prod_wo_range4010w(0) <= lsb_prod_wo(29);
	wire_man_prod_w_lsb_prod_wo_range4172w(0) <= lsb_prod_wo(2);
	wire_man_prod_w_lsb_prod_wo_range4004w(0) <= lsb_prod_wo(30);
	wire_man_prod_w_lsb_prod_wo_range3998w(0) <= lsb_prod_wo(31);
	wire_man_prod_w_lsb_prod_wo_range3992w(0) <= lsb_prod_wo(32);
	wire_man_prod_w_lsb_prod_wo_range3986w(0) <= lsb_prod_wo(33);
	wire_man_prod_w_lsb_prod_wo_range3980w(0) <= lsb_prod_wo(34);
	wire_man_prod_w_lsb_prod_wo_range3974w(0) <= lsb_prod_wo(35);
	wire_man_prod_w_lsb_prod_wo_range3968w(0) <= lsb_prod_wo(36);
	wire_man_prod_w_lsb_prod_wo_range3962w(0) <= lsb_prod_wo(37);
	wire_man_prod_w_lsb_prod_wo_range3956w(0) <= lsb_prod_wo(38);
	wire_man_prod_w_lsb_prod_wo_range3950w(0) <= lsb_prod_wo(39);
	wire_man_prod_w_lsb_prod_wo_range4166w(0) <= lsb_prod_wo(3);
	wire_man_prod_w_lsb_prod_wo_range3944w(0) <= lsb_prod_wo(40);
	wire_man_prod_w_lsb_prod_wo_range3938w(0) <= lsb_prod_wo(41);
	wire_man_prod_w_lsb_prod_wo_range3932w(0) <= lsb_prod_wo(42);
	wire_man_prod_w_lsb_prod_wo_range3926w(0) <= lsb_prod_wo(43);
	wire_man_prod_w_lsb_prod_wo_range3920w(0) <= lsb_prod_wo(44);
	wire_man_prod_w_lsb_prod_wo_range3914w(0) <= lsb_prod_wo(45);
	wire_man_prod_w_lsb_prod_wo_range3908w(0) <= lsb_prod_wo(46);
	wire_man_prod_w_lsb_prod_wo_range3902w(0) <= lsb_prod_wo(47);
	wire_man_prod_w_lsb_prod_wo_range3896w(0) <= lsb_prod_wo(48);
	wire_man_prod_w_lsb_prod_wo_range3890w(0) <= lsb_prod_wo(49);
	wire_man_prod_w_lsb_prod_wo_range4160w(0) <= lsb_prod_wo(4);
	wire_man_prod_w_lsb_prod_wo_range3884w(0) <= lsb_prod_wo(50);
	wire_man_prod_w_lsb_prod_wo_range3878w(0) <= lsb_prod_wo(51);
	wire_man_prod_w_lsb_prod_wo_range3872w(0) <= lsb_prod_wo(52);
	wire_man_prod_w_lsb_prod_wo_range3866w(0) <= lsb_prod_wo(53);
	wire_man_prod_w_lsb_prod_wo_range3860w(0) <= lsb_prod_wo(54);
	wire_man_prod_w_lsb_prod_wo_range3854w(0) <= lsb_prod_wo(55);
	wire_man_prod_w_lsb_prod_wo_range3848w(0) <= lsb_prod_wo(56);
	wire_man_prod_w_lsb_prod_wo_range3842w(0) <= lsb_prod_wo(57);
	wire_man_prod_w_lsb_prod_wo_range3836w(0) <= lsb_prod_wo(58);
	wire_man_prod_w_lsb_prod_wo_range3830w(0) <= lsb_prod_wo(59);
	wire_man_prod_w_lsb_prod_wo_range4154w(0) <= lsb_prod_wo(5);
	wire_man_prod_w_lsb_prod_wo_range4148w(0) <= lsb_prod_wo(6);
	wire_man_prod_w_lsb_prod_wo_range4142w(0) <= lsb_prod_wo(7);
	wire_man_prod_w_lsb_prod_wo_range4136w(0) <= lsb_prod_wo(8);
	wire_man_prod_w_lsb_prod_wo_range4130w(0) <= lsb_prod_wo(9);
	wire_man_prod_w_msb_prod_wo_range4181w(0) <= msb_prod_wo(0);
	wire_man_prod_w_msb_prod_wo_range4121w(0) <= msb_prod_wo(10);
	wire_man_prod_w_msb_prod_wo_range4115w(0) <= msb_prod_wo(11);
	wire_man_prod_w_msb_prod_wo_range4109w(0) <= msb_prod_wo(12);
	wire_man_prod_w_msb_prod_wo_range4103w(0) <= msb_prod_wo(13);
	wire_man_prod_w_msb_prod_wo_range4097w(0) <= msb_prod_wo(14);
	wire_man_prod_w_msb_prod_wo_range4091w(0) <= msb_prod_wo(15);
	wire_man_prod_w_msb_prod_wo_range4085w(0) <= msb_prod_wo(16);
	wire_man_prod_w_msb_prod_wo_range4079w(0) <= msb_prod_wo(17);
	wire_man_prod_w_msb_prod_wo_range4073w(0) <= msb_prod_wo(18);
	wire_man_prod_w_msb_prod_wo_range4067w(0) <= msb_prod_wo(19);
	wire_man_prod_w_msb_prod_wo_range4175w(0) <= msb_prod_wo(1);
	wire_man_prod_w_msb_prod_wo_range4061w(0) <= msb_prod_wo(20);
	wire_man_prod_w_msb_prod_wo_range4055w(0) <= msb_prod_wo(21);
	wire_man_prod_w_msb_prod_wo_range4049w(0) <= msb_prod_wo(22);
	wire_man_prod_w_msb_prod_wo_range4043w(0) <= msb_prod_wo(23);
	wire_man_prod_w_msb_prod_wo_range4037w(0) <= msb_prod_wo(24);
	wire_man_prod_w_msb_prod_wo_range4031w(0) <= msb_prod_wo(25);
	wire_man_prod_w_msb_prod_wo_range4025w(0) <= msb_prod_wo(26);
	wire_man_prod_w_msb_prod_wo_range4019w(0) <= msb_prod_wo(27);
	wire_man_prod_w_msb_prod_wo_range4013w(0) <= msb_prod_wo(28);
	wire_man_prod_w_msb_prod_wo_range4007w(0) <= msb_prod_wo(29);
	wire_man_prod_w_msb_prod_wo_range4169w(0) <= msb_prod_wo(2);
	wire_man_prod_w_msb_prod_wo_range4001w(0) <= msb_prod_wo(30);
	wire_man_prod_w_msb_prod_wo_range3995w(0) <= msb_prod_wo(31);
	wire_man_prod_w_msb_prod_wo_range3989w(0) <= msb_prod_wo(32);
	wire_man_prod_w_msb_prod_wo_range3983w(0) <= msb_prod_wo(33);
	wire_man_prod_w_msb_prod_wo_range3977w(0) <= msb_prod_wo(34);
	wire_man_prod_w_msb_prod_wo_range3971w(0) <= msb_prod_wo(35);
	wire_man_prod_w_msb_prod_wo_range3965w(0) <= msb_prod_wo(36);
	wire_man_prod_w_msb_prod_wo_range3959w(0) <= msb_prod_wo(37);
	wire_man_prod_w_msb_prod_wo_range3953w(0) <= msb_prod_wo(38);
	wire_man_prod_w_msb_prod_wo_range3947w(0) <= msb_prod_wo(39);
	wire_man_prod_w_msb_prod_wo_range4163w(0) <= msb_prod_wo(3);
	wire_man_prod_w_msb_prod_wo_range3941w(0) <= msb_prod_wo(40);
	wire_man_prod_w_msb_prod_wo_range3935w(0) <= msb_prod_wo(41);
	wire_man_prod_w_msb_prod_wo_range3929w(0) <= msb_prod_wo(42);
	wire_man_prod_w_msb_prod_wo_range3923w(0) <= msb_prod_wo(43);
	wire_man_prod_w_msb_prod_wo_range3917w(0) <= msb_prod_wo(44);
	wire_man_prod_w_msb_prod_wo_range3911w(0) <= msb_prod_wo(45);
	wire_man_prod_w_msb_prod_wo_range3905w(0) <= msb_prod_wo(46);
	wire_man_prod_w_msb_prod_wo_range3899w(0) <= msb_prod_wo(47);
	wire_man_prod_w_msb_prod_wo_range3893w(0) <= msb_prod_wo(48);
	wire_man_prod_w_msb_prod_wo_range3887w(0) <= msb_prod_wo(49);
	wire_man_prod_w_msb_prod_wo_range4157w(0) <= msb_prod_wo(4);
	wire_man_prod_w_msb_prod_wo_range3881w(0) <= msb_prod_wo(50);
	wire_man_prod_w_msb_prod_wo_range3875w(0) <= msb_prod_wo(51);
	wire_man_prod_w_msb_prod_wo_range3869w(0) <= msb_prod_wo(52);
	wire_man_prod_w_msb_prod_wo_range3863w(0) <= msb_prod_wo(53);
	wire_man_prod_w_msb_prod_wo_range3857w(0) <= msb_prod_wo(54);
	wire_man_prod_w_msb_prod_wo_range3851w(0) <= msb_prod_wo(55);
	wire_man_prod_w_msb_prod_wo_range3845w(0) <= msb_prod_wo(56);
	wire_man_prod_w_msb_prod_wo_range3839w(0) <= msb_prod_wo(57);
	wire_man_prod_w_msb_prod_wo_range3833w(0) <= msb_prod_wo(58);
	wire_man_prod_w_msb_prod_wo_range3827w(0) <= msb_prod_wo(59);
	wire_man_prod_w_msb_prod_wo_range4151w(0) <= msb_prod_wo(5);
	wire_man_prod_w_msb_prod_wo_range4145w(0) <= msb_prod_wo(6);
	wire_man_prod_w_msb_prod_wo_range4139w(0) <= msb_prod_wo(7);
	wire_man_prod_w_msb_prod_wo_range4133w(0) <= msb_prod_wo(8);
	wire_man_prod_w_msb_prod_wo_range4127w(0) <= msb_prod_wo(9);
	wire_man_prod_w_neg_lsb_range4186w(0) <= neg_lsb(0);
	wire_man_prod_w_neg_lsb_range4126w(0) <= neg_lsb(10);
	wire_man_prod_w_neg_lsb_range4120w(0) <= neg_lsb(11);
	wire_man_prod_w_neg_lsb_range4114w(0) <= neg_lsb(12);
	wire_man_prod_w_neg_lsb_range4108w(0) <= neg_lsb(13);
	wire_man_prod_w_neg_lsb_range4102w(0) <= neg_lsb(14);
	wire_man_prod_w_neg_lsb_range4096w(0) <= neg_lsb(15);
	wire_man_prod_w_neg_lsb_range4090w(0) <= neg_lsb(16);
	wire_man_prod_w_neg_lsb_range4084w(0) <= neg_lsb(17);
	wire_man_prod_w_neg_lsb_range4078w(0) <= neg_lsb(18);
	wire_man_prod_w_neg_lsb_range4072w(0) <= neg_lsb(19);
	wire_man_prod_w_neg_lsb_range4180w(0) <= neg_lsb(1);
	wire_man_prod_w_neg_lsb_range4066w(0) <= neg_lsb(20);
	wire_man_prod_w_neg_lsb_range4060w(0) <= neg_lsb(21);
	wire_man_prod_w_neg_lsb_range4054w(0) <= neg_lsb(22);
	wire_man_prod_w_neg_lsb_range4048w(0) <= neg_lsb(23);
	wire_man_prod_w_neg_lsb_range4042w(0) <= neg_lsb(24);
	wire_man_prod_w_neg_lsb_range4036w(0) <= neg_lsb(25);
	wire_man_prod_w_neg_lsb_range4030w(0) <= neg_lsb(26);
	wire_man_prod_w_neg_lsb_range4024w(0) <= neg_lsb(27);
	wire_man_prod_w_neg_lsb_range4018w(0) <= neg_lsb(28);
	wire_man_prod_w_neg_lsb_range4012w(0) <= neg_lsb(29);
	wire_man_prod_w_neg_lsb_range4174w(0) <= neg_lsb(2);
	wire_man_prod_w_neg_lsb_range4006w(0) <= neg_lsb(30);
	wire_man_prod_w_neg_lsb_range4000w(0) <= neg_lsb(31);
	wire_man_prod_w_neg_lsb_range3994w(0) <= neg_lsb(32);
	wire_man_prod_w_neg_lsb_range3988w(0) <= neg_lsb(33);
	wire_man_prod_w_neg_lsb_range3982w(0) <= neg_lsb(34);
	wire_man_prod_w_neg_lsb_range3976w(0) <= neg_lsb(35);
	wire_man_prod_w_neg_lsb_range3970w(0) <= neg_lsb(36);
	wire_man_prod_w_neg_lsb_range3964w(0) <= neg_lsb(37);
	wire_man_prod_w_neg_lsb_range3958w(0) <= neg_lsb(38);
	wire_man_prod_w_neg_lsb_range3952w(0) <= neg_lsb(39);
	wire_man_prod_w_neg_lsb_range4168w(0) <= neg_lsb(3);
	wire_man_prod_w_neg_lsb_range3946w(0) <= neg_lsb(40);
	wire_man_prod_w_neg_lsb_range3940w(0) <= neg_lsb(41);
	wire_man_prod_w_neg_lsb_range3934w(0) <= neg_lsb(42);
	wire_man_prod_w_neg_lsb_range3928w(0) <= neg_lsb(43);
	wire_man_prod_w_neg_lsb_range3922w(0) <= neg_lsb(44);
	wire_man_prod_w_neg_lsb_range3916w(0) <= neg_lsb(45);
	wire_man_prod_w_neg_lsb_range3910w(0) <= neg_lsb(46);
	wire_man_prod_w_neg_lsb_range3904w(0) <= neg_lsb(47);
	wire_man_prod_w_neg_lsb_range3898w(0) <= neg_lsb(48);
	wire_man_prod_w_neg_lsb_range3892w(0) <= neg_lsb(49);
	wire_man_prod_w_neg_lsb_range4162w(0) <= neg_lsb(4);
	wire_man_prod_w_neg_lsb_range3886w(0) <= neg_lsb(50);
	wire_man_prod_w_neg_lsb_range3880w(0) <= neg_lsb(51);
	wire_man_prod_w_neg_lsb_range3874w(0) <= neg_lsb(52);
	wire_man_prod_w_neg_lsb_range3868w(0) <= neg_lsb(53);
	wire_man_prod_w_neg_lsb_range3862w(0) <= neg_lsb(54);
	wire_man_prod_w_neg_lsb_range3856w(0) <= neg_lsb(55);
	wire_man_prod_w_neg_lsb_range3850w(0) <= neg_lsb(56);
	wire_man_prod_w_neg_lsb_range3844w(0) <= neg_lsb(57);
	wire_man_prod_w_neg_lsb_range3838w(0) <= neg_lsb(58);
	wire_man_prod_w_neg_lsb_range3832w(0) <= neg_lsb(59);
	wire_man_prod_w_neg_lsb_range4156w(0) <= neg_lsb(5);
	wire_man_prod_w_neg_lsb_range3825w(0) <= neg_lsb(60);
	wire_man_prod_w_neg_lsb_range3821w(0) <= neg_lsb(61);
	wire_man_prod_w_neg_lsb_range3817w(0) <= neg_lsb(62);
	wire_man_prod_w_neg_lsb_range3813w(0) <= neg_lsb(63);
	wire_man_prod_w_neg_lsb_range3809w(0) <= neg_lsb(64);
	wire_man_prod_w_neg_lsb_range3805w(0) <= neg_lsb(65);
	wire_man_prod_w_neg_lsb_range3801w(0) <= neg_lsb(66);
	wire_man_prod_w_neg_lsb_range3797w(0) <= neg_lsb(67);
	wire_man_prod_w_neg_lsb_range3793w(0) <= neg_lsb(68);
	wire_man_prod_w_neg_lsb_range3789w(0) <= neg_lsb(69);
	wire_man_prod_w_neg_lsb_range4150w(0) <= neg_lsb(6);
	wire_man_prod_w_neg_lsb_range3785w(0) <= neg_lsb(70);
	wire_man_prod_w_neg_lsb_range3781w(0) <= neg_lsb(71);
	wire_man_prod_w_neg_lsb_range3777w(0) <= neg_lsb(72);
	wire_man_prod_w_neg_lsb_range3773w(0) <= neg_lsb(73);
	wire_man_prod_w_neg_lsb_range3769w(0) <= neg_lsb(74);
	wire_man_prod_w_neg_lsb_range3765w(0) <= neg_lsb(75);
	wire_man_prod_w_neg_lsb_range3761w(0) <= neg_lsb(76);
	wire_man_prod_w_neg_lsb_range3757w(0) <= neg_lsb(77);
	wire_man_prod_w_neg_lsb_range3753w(0) <= neg_lsb(78);
	wire_man_prod_w_neg_lsb_range3749w(0) <= neg_lsb(79);
	wire_man_prod_w_neg_lsb_range4144w(0) <= neg_lsb(7);
	wire_man_prod_w_neg_lsb_range3745w(0) <= neg_lsb(80);
	wire_man_prod_w_neg_lsb_range3741w(0) <= neg_lsb(81);
	wire_man_prod_w_neg_lsb_range3737w(0) <= neg_lsb(82);
	wire_man_prod_w_neg_lsb_range3733w(0) <= neg_lsb(83);
	wire_man_prod_w_neg_lsb_range3729w(0) <= neg_lsb(84);
	wire_man_prod_w_neg_lsb_range3725w(0) <= neg_lsb(85);
	wire_man_prod_w_neg_lsb_range3721w(0) <= neg_lsb(86);
	wire_man_prod_w_neg_lsb_range3717w(0) <= neg_lsb(87);
	wire_man_prod_w_neg_lsb_range3713w(0) <= neg_lsb(88);
	wire_man_prod_w_neg_lsb_range3708w(0) <= neg_lsb(89);
	wire_man_prod_w_neg_lsb_range4138w(0) <= neg_lsb(8);
	wire_man_prod_w_neg_lsb_range4132w(0) <= neg_lsb(9);
	wire_man_prod_w_neg_msb_range4183w(0) <= neg_msb(0);
	wire_man_prod_w_neg_msb_range4123w(0) <= neg_msb(10);
	wire_man_prod_w_neg_msb_range4117w(0) <= neg_msb(11);
	wire_man_prod_w_neg_msb_range4111w(0) <= neg_msb(12);
	wire_man_prod_w_neg_msb_range4105w(0) <= neg_msb(13);
	wire_man_prod_w_neg_msb_range4099w(0) <= neg_msb(14);
	wire_man_prod_w_neg_msb_range4093w(0) <= neg_msb(15);
	wire_man_prod_w_neg_msb_range4087w(0) <= neg_msb(16);
	wire_man_prod_w_neg_msb_range4081w(0) <= neg_msb(17);
	wire_man_prod_w_neg_msb_range4075w(0) <= neg_msb(18);
	wire_man_prod_w_neg_msb_range4069w(0) <= neg_msb(19);
	wire_man_prod_w_neg_msb_range4177w(0) <= neg_msb(1);
	wire_man_prod_w_neg_msb_range4063w(0) <= neg_msb(20);
	wire_man_prod_w_neg_msb_range4057w(0) <= neg_msb(21);
	wire_man_prod_w_neg_msb_range4051w(0) <= neg_msb(22);
	wire_man_prod_w_neg_msb_range4045w(0) <= neg_msb(23);
	wire_man_prod_w_neg_msb_range4039w(0) <= neg_msb(24);
	wire_man_prod_w_neg_msb_range4033w(0) <= neg_msb(25);
	wire_man_prod_w_neg_msb_range4027w(0) <= neg_msb(26);
	wire_man_prod_w_neg_msb_range4021w(0) <= neg_msb(27);
	wire_man_prod_w_neg_msb_range4015w(0) <= neg_msb(28);
	wire_man_prod_w_neg_msb_range4009w(0) <= neg_msb(29);
	wire_man_prod_w_neg_msb_range4171w(0) <= neg_msb(2);
	wire_man_prod_w_neg_msb_range4003w(0) <= neg_msb(30);
	wire_man_prod_w_neg_msb_range3997w(0) <= neg_msb(31);
	wire_man_prod_w_neg_msb_range3991w(0) <= neg_msb(32);
	wire_man_prod_w_neg_msb_range3985w(0) <= neg_msb(33);
	wire_man_prod_w_neg_msb_range3979w(0) <= neg_msb(34);
	wire_man_prod_w_neg_msb_range3973w(0) <= neg_msb(35);
	wire_man_prod_w_neg_msb_range3967w(0) <= neg_msb(36);
	wire_man_prod_w_neg_msb_range3961w(0) <= neg_msb(37);
	wire_man_prod_w_neg_msb_range3955w(0) <= neg_msb(38);
	wire_man_prod_w_neg_msb_range3949w(0) <= neg_msb(39);
	wire_man_prod_w_neg_msb_range4165w(0) <= neg_msb(3);
	wire_man_prod_w_neg_msb_range3943w(0) <= neg_msb(40);
	wire_man_prod_w_neg_msb_range3937w(0) <= neg_msb(41);
	wire_man_prod_w_neg_msb_range3931w(0) <= neg_msb(42);
	wire_man_prod_w_neg_msb_range3925w(0) <= neg_msb(43);
	wire_man_prod_w_neg_msb_range3919w(0) <= neg_msb(44);
	wire_man_prod_w_neg_msb_range3913w(0) <= neg_msb(45);
	wire_man_prod_w_neg_msb_range3907w(0) <= neg_msb(46);
	wire_man_prod_w_neg_msb_range3901w(0) <= neg_msb(47);
	wire_man_prod_w_neg_msb_range3895w(0) <= neg_msb(48);
	wire_man_prod_w_neg_msb_range3889w(0) <= neg_msb(49);
	wire_man_prod_w_neg_msb_range4159w(0) <= neg_msb(4);
	wire_man_prod_w_neg_msb_range3883w(0) <= neg_msb(50);
	wire_man_prod_w_neg_msb_range3877w(0) <= neg_msb(51);
	wire_man_prod_w_neg_msb_range3871w(0) <= neg_msb(52);
	wire_man_prod_w_neg_msb_range3865w(0) <= neg_msb(53);
	wire_man_prod_w_neg_msb_range3859w(0) <= neg_msb(54);
	wire_man_prod_w_neg_msb_range3853w(0) <= neg_msb(55);
	wire_man_prod_w_neg_msb_range3847w(0) <= neg_msb(56);
	wire_man_prod_w_neg_msb_range3841w(0) <= neg_msb(57);
	wire_man_prod_w_neg_msb_range3835w(0) <= neg_msb(58);
	wire_man_prod_w_neg_msb_range3829w(0) <= neg_msb(59);
	wire_man_prod_w_neg_msb_range4153w(0) <= neg_msb(5);
	wire_man_prod_w_neg_msb_range3823w(0) <= neg_msb(60);
	wire_man_prod_w_neg_msb_range3819w(0) <= neg_msb(61);
	wire_man_prod_w_neg_msb_range3815w(0) <= neg_msb(62);
	wire_man_prod_w_neg_msb_range3811w(0) <= neg_msb(63);
	wire_man_prod_w_neg_msb_range3807w(0) <= neg_msb(64);
	wire_man_prod_w_neg_msb_range3803w(0) <= neg_msb(65);
	wire_man_prod_w_neg_msb_range3799w(0) <= neg_msb(66);
	wire_man_prod_w_neg_msb_range3795w(0) <= neg_msb(67);
	wire_man_prod_w_neg_msb_range3791w(0) <= neg_msb(68);
	wire_man_prod_w_neg_msb_range3787w(0) <= neg_msb(69);
	wire_man_prod_w_neg_msb_range4147w(0) <= neg_msb(6);
	wire_man_prod_w_neg_msb_range3783w(0) <= neg_msb(70);
	wire_man_prod_w_neg_msb_range3779w(0) <= neg_msb(71);
	wire_man_prod_w_neg_msb_range3775w(0) <= neg_msb(72);
	wire_man_prod_w_neg_msb_range3771w(0) <= neg_msb(73);
	wire_man_prod_w_neg_msb_range3767w(0) <= neg_msb(74);
	wire_man_prod_w_neg_msb_range3763w(0) <= neg_msb(75);
	wire_man_prod_w_neg_msb_range3759w(0) <= neg_msb(76);
	wire_man_prod_w_neg_msb_range3755w(0) <= neg_msb(77);
	wire_man_prod_w_neg_msb_range3751w(0) <= neg_msb(78);
	wire_man_prod_w_neg_msb_range3747w(0) <= neg_msb(79);
	wire_man_prod_w_neg_msb_range4141w(0) <= neg_msb(7);
	wire_man_prod_w_neg_msb_range3743w(0) <= neg_msb(80);
	wire_man_prod_w_neg_msb_range3739w(0) <= neg_msb(81);
	wire_man_prod_w_neg_msb_range3735w(0) <= neg_msb(82);
	wire_man_prod_w_neg_msb_range3731w(0) <= neg_msb(83);
	wire_man_prod_w_neg_msb_range3727w(0) <= neg_msb(84);
	wire_man_prod_w_neg_msb_range3723w(0) <= neg_msb(85);
	wire_man_prod_w_neg_msb_range3719w(0) <= neg_msb(86);
	wire_man_prod_w_neg_msb_range3715w(0) <= neg_msb(87);
	wire_man_prod_w_neg_msb_range3711w(0) <= neg_msb(88);
	wire_man_prod_w_neg_msb_range3705w(0) <= neg_msb(89);
	wire_man_prod_w_neg_msb_range4135w(0) <= neg_msb(8);
	wire_man_prod_w_neg_msb_range4129w(0) <= neg_msb(9);
	wire_man_prod_w_sum_one_range4190w(0) <= sum_one(0);
	wire_man_prod_w_sum_one_range4292w(0) <= sum_one(10);
	wire_man_prod_w_sum_one_range4302w(0) <= sum_one(11);
	wire_man_prod_w_sum_one_range4312w(0) <= sum_one(12);
	wire_man_prod_w_sum_one_range4322w(0) <= sum_one(13);
	wire_man_prod_w_sum_one_range4332w(0) <= sum_one(14);
	wire_man_prod_w_sum_one_range4342w(0) <= sum_one(15);
	wire_man_prod_w_sum_one_range4352w(0) <= sum_one(16);
	wire_man_prod_w_sum_one_range4362w(0) <= sum_one(17);
	wire_man_prod_w_sum_one_range4372w(0) <= sum_one(18);
	wire_man_prod_w_sum_one_range4382w(0) <= sum_one(19);
	wire_man_prod_w_sum_one_range4202w(0) <= sum_one(1);
	wire_man_prod_w_sum_one_range4392w(0) <= sum_one(20);
	wire_man_prod_w_sum_one_range4402w(0) <= sum_one(21);
	wire_man_prod_w_sum_one_range4412w(0) <= sum_one(22);
	wire_man_prod_w_sum_one_range4422w(0) <= sum_one(23);
	wire_man_prod_w_sum_one_range4432w(0) <= sum_one(24);
	wire_man_prod_w_sum_one_range4442w(0) <= sum_one(25);
	wire_man_prod_w_sum_one_range4452w(0) <= sum_one(26);
	wire_man_prod_w_sum_one_range4462w(0) <= sum_one(27);
	wire_man_prod_w_sum_one_range4472w(0) <= sum_one(28);
	wire_man_prod_w_sum_one_range4482w(0) <= sum_one(29);
	wire_man_prod_w_sum_one_range4212w(0) <= sum_one(2);
	wire_man_prod_w_sum_one_range4492w(0) <= sum_one(30);
	wire_man_prod_w_sum_one_range4502w(0) <= sum_one(31);
	wire_man_prod_w_sum_one_range4512w(0) <= sum_one(32);
	wire_man_prod_w_sum_one_range4522w(0) <= sum_one(33);
	wire_man_prod_w_sum_one_range4532w(0) <= sum_one(34);
	wire_man_prod_w_sum_one_range4542w(0) <= sum_one(35);
	wire_man_prod_w_sum_one_range4552w(0) <= sum_one(36);
	wire_man_prod_w_sum_one_range4562w(0) <= sum_one(37);
	wire_man_prod_w_sum_one_range4572w(0) <= sum_one(38);
	wire_man_prod_w_sum_one_range4582w(0) <= sum_one(39);
	wire_man_prod_w_sum_one_range4222w(0) <= sum_one(3);
	wire_man_prod_w_sum_one_range4592w(0) <= sum_one(40);
	wire_man_prod_w_sum_one_range4602w(0) <= sum_one(41);
	wire_man_prod_w_sum_one_range4612w(0) <= sum_one(42);
	wire_man_prod_w_sum_one_range4622w(0) <= sum_one(43);
	wire_man_prod_w_sum_one_range4632w(0) <= sum_one(44);
	wire_man_prod_w_sum_one_range4642w(0) <= sum_one(45);
	wire_man_prod_w_sum_one_range4652w(0) <= sum_one(46);
	wire_man_prod_w_sum_one_range4662w(0) <= sum_one(47);
	wire_man_prod_w_sum_one_range4672w(0) <= sum_one(48);
	wire_man_prod_w_sum_one_range4682w(0) <= sum_one(49);
	wire_man_prod_w_sum_one_range4232w(0) <= sum_one(4);
	wire_man_prod_w_sum_one_range4692w(0) <= sum_one(50);
	wire_man_prod_w_sum_one_range4702w(0) <= sum_one(51);
	wire_man_prod_w_sum_one_range4712w(0) <= sum_one(52);
	wire_man_prod_w_sum_one_range4722w(0) <= sum_one(53);
	wire_man_prod_w_sum_one_range4732w(0) <= sum_one(54);
	wire_man_prod_w_sum_one_range4742w(0) <= sum_one(55);
	wire_man_prod_w_sum_one_range4752w(0) <= sum_one(56);
	wire_man_prod_w_sum_one_range4762w(0) <= sum_one(57);
	wire_man_prod_w_sum_one_range4772w(0) <= sum_one(58);
	wire_man_prod_w_sum_one_range4782w(0) <= sum_one(59);
	wire_man_prod_w_sum_one_range4242w(0) <= sum_one(5);
	wire_man_prod_w_sum_one_range4792w(0) <= sum_one(60);
	wire_man_prod_w_sum_one_range4802w(0) <= sum_one(61);
	wire_man_prod_w_sum_one_range4812w(0) <= sum_one(62);
	wire_man_prod_w_sum_one_range4822w(0) <= sum_one(63);
	wire_man_prod_w_sum_one_range4832w(0) <= sum_one(64);
	wire_man_prod_w_sum_one_range4842w(0) <= sum_one(65);
	wire_man_prod_w_sum_one_range4852w(0) <= sum_one(66);
	wire_man_prod_w_sum_one_range4862w(0) <= sum_one(67);
	wire_man_prod_w_sum_one_range4872w(0) <= sum_one(68);
	wire_man_prod_w_sum_one_range4882w(0) <= sum_one(69);
	wire_man_prod_w_sum_one_range4252w(0) <= sum_one(6);
	wire_man_prod_w_sum_one_range4892w(0) <= sum_one(70);
	wire_man_prod_w_sum_one_range4902w(0) <= sum_one(71);
	wire_man_prod_w_sum_one_range4912w(0) <= sum_one(72);
	wire_man_prod_w_sum_one_range4922w(0) <= sum_one(73);
	wire_man_prod_w_sum_one_range4932w(0) <= sum_one(74);
	wire_man_prod_w_sum_one_range4942w(0) <= sum_one(75);
	wire_man_prod_w_sum_one_range4952w(0) <= sum_one(76);
	wire_man_prod_w_sum_one_range4962w(0) <= sum_one(77);
	wire_man_prod_w_sum_one_range4972w(0) <= sum_one(78);
	wire_man_prod_w_sum_one_range4982w(0) <= sum_one(79);
	wire_man_prod_w_sum_one_range4262w(0) <= sum_one(7);
	wire_man_prod_w_sum_one_range4992w(0) <= sum_one(80);
	wire_man_prod_w_sum_one_range5002w(0) <= sum_one(81);
	wire_man_prod_w_sum_one_range5012w(0) <= sum_one(82);
	wire_man_prod_w_sum_one_range5022w(0) <= sum_one(83);
	wire_man_prod_w_sum_one_range5032w(0) <= sum_one(84);
	wire_man_prod_w_sum_one_range5042w(0) <= sum_one(85);
	wire_man_prod_w_sum_one_range5052w(0) <= sum_one(86);
	wire_man_prod_w_sum_one_range5062w(0) <= sum_one(87);
	wire_man_prod_w_sum_one_range5072w(0) <= sum_one(88);
	wire_man_prod_w_sum_one_range5082w(0) <= sum_one(89);
	wire_man_prod_w_sum_one_range4272w(0) <= sum_one(8);
	wire_man_prod_w_sum_one_range4282w(0) <= sum_one(9);
	wire_man_prod_w_vector1_range5094w(0) <= vector1(0);
	wire_man_prod_w_vector1_range5206w(0) <= vector1(10);
	wire_man_prod_w_vector1_range5217w(0) <= vector1(11);
	wire_man_prod_w_vector1_range5228w(0) <= vector1(12);
	wire_man_prod_w_vector1_range5239w(0) <= vector1(13);
	wire_man_prod_w_vector1_range5250w(0) <= vector1(14);
	wire_man_prod_w_vector1_range5261w(0) <= vector1(15);
	wire_man_prod_w_vector1_range5272w(0) <= vector1(16);
	wire_man_prod_w_vector1_range5283w(0) <= vector1(17);
	wire_man_prod_w_vector1_range5294w(0) <= vector1(18);
	wire_man_prod_w_vector1_range5305w(0) <= vector1(19);
	wire_man_prod_w_vector1_range5107w(0) <= vector1(1);
	wire_man_prod_w_vector1_range5316w(0) <= vector1(20);
	wire_man_prod_w_vector1_range5327w(0) <= vector1(21);
	wire_man_prod_w_vector1_range5338w(0) <= vector1(22);
	wire_man_prod_w_vector1_range5349w(0) <= vector1(23);
	wire_man_prod_w_vector1_range5360w(0) <= vector1(24);
	wire_man_prod_w_vector1_range5371w(0) <= vector1(25);
	wire_man_prod_w_vector1_range5382w(0) <= vector1(26);
	wire_man_prod_w_vector1_range5393w(0) <= vector1(27);
	wire_man_prod_w_vector1_range5404w(0) <= vector1(28);
	wire_man_prod_w_vector1_range5415w(0) <= vector1(29);
	wire_man_prod_w_vector1_range5118w(0) <= vector1(2);
	wire_man_prod_w_vector1_range5426w(0) <= vector1(30);
	wire_man_prod_w_vector1_range5437w(0) <= vector1(31);
	wire_man_prod_w_vector1_range5448w(0) <= vector1(32);
	wire_man_prod_w_vector1_range5459w(0) <= vector1(33);
	wire_man_prod_w_vector1_range5470w(0) <= vector1(34);
	wire_man_prod_w_vector1_range5481w(0) <= vector1(35);
	wire_man_prod_w_vector1_range5492w(0) <= vector1(36);
	wire_man_prod_w_vector1_range5503w(0) <= vector1(37);
	wire_man_prod_w_vector1_range5514w(0) <= vector1(38);
	wire_man_prod_w_vector1_range5525w(0) <= vector1(39);
	wire_man_prod_w_vector1_range5129w(0) <= vector1(3);
	wire_man_prod_w_vector1_range5536w(0) <= vector1(40);
	wire_man_prod_w_vector1_range5547w(0) <= vector1(41);
	wire_man_prod_w_vector1_range5558w(0) <= vector1(42);
	wire_man_prod_w_vector1_range5569w(0) <= vector1(43);
	wire_man_prod_w_vector1_range5580w(0) <= vector1(44);
	wire_man_prod_w_vector1_range5591w(0) <= vector1(45);
	wire_man_prod_w_vector1_range5602w(0) <= vector1(46);
	wire_man_prod_w_vector1_range5613w(0) <= vector1(47);
	wire_man_prod_w_vector1_range5624w(0) <= vector1(48);
	wire_man_prod_w_vector1_range5635w(0) <= vector1(49);
	wire_man_prod_w_vector1_range5140w(0) <= vector1(4);
	wire_man_prod_w_vector1_range5646w(0) <= vector1(50);
	wire_man_prod_w_vector1_range5657w(0) <= vector1(51);
	wire_man_prod_w_vector1_range5668w(0) <= vector1(52);
	wire_man_prod_w_vector1_range5679w(0) <= vector1(53);
	wire_man_prod_w_vector1_range5690w(0) <= vector1(54);
	wire_man_prod_w_vector1_range5701w(0) <= vector1(55);
	wire_man_prod_w_vector1_range5712w(0) <= vector1(56);
	wire_man_prod_w_vector1_range5723w(0) <= vector1(57);
	wire_man_prod_w_vector1_range5734w(0) <= vector1(58);
	wire_man_prod_w_vector1_range5745w(0) <= vector1(59);
	wire_man_prod_w_vector1_range5151w(0) <= vector1(5);
	wire_man_prod_w_vector1_range5756w(0) <= vector1(60);
	wire_man_prod_w_vector1_range5767w(0) <= vector1(61);
	wire_man_prod_w_vector1_range5778w(0) <= vector1(62);
	wire_man_prod_w_vector1_range5789w(0) <= vector1(63);
	wire_man_prod_w_vector1_range5800w(0) <= vector1(64);
	wire_man_prod_w_vector1_range5811w(0) <= vector1(65);
	wire_man_prod_w_vector1_range5822w(0) <= vector1(66);
	wire_man_prod_w_vector1_range5833w(0) <= vector1(67);
	wire_man_prod_w_vector1_range5844w(0) <= vector1(68);
	wire_man_prod_w_vector1_range5855w(0) <= vector1(69);
	wire_man_prod_w_vector1_range5162w(0) <= vector1(6);
	wire_man_prod_w_vector1_range5866w(0) <= vector1(70);
	wire_man_prod_w_vector1_range5877w(0) <= vector1(71);
	wire_man_prod_w_vector1_range5888w(0) <= vector1(72);
	wire_man_prod_w_vector1_range5899w(0) <= vector1(73);
	wire_man_prod_w_vector1_range5910w(0) <= vector1(74);
	wire_man_prod_w_vector1_range5921w(0) <= vector1(75);
	wire_man_prod_w_vector1_range5932w(0) <= vector1(76);
	wire_man_prod_w_vector1_range5943w(0) <= vector1(77);
	wire_man_prod_w_vector1_range5954w(0) <= vector1(78);
	wire_man_prod_w_vector1_range5965w(0) <= vector1(79);
	wire_man_prod_w_vector1_range5173w(0) <= vector1(7);
	wire_man_prod_w_vector1_range5976w(0) <= vector1(80);
	wire_man_prod_w_vector1_range5987w(0) <= vector1(81);
	wire_man_prod_w_vector1_range5998w(0) <= vector1(82);
	wire_man_prod_w_vector1_range6009w(0) <= vector1(83);
	wire_man_prod_w_vector1_range6020w(0) <= vector1(84);
	wire_man_prod_w_vector1_range6031w(0) <= vector1(85);
	wire_man_prod_w_vector1_range6042w(0) <= vector1(86);
	wire_man_prod_w_vector1_range6053w(0) <= vector1(87);
	wire_man_prod_w_vector1_range6064w(0) <= vector1(88);
	wire_man_prod_w_vector1_range6075w(0) <= vector1(89);
	wire_man_prod_w_vector1_range5184w(0) <= vector1(8);
	wire_man_prod_w_vector1_range5195w(0) <= vector1(9);
	wire_man_prod_w_vector2_range4187w(0) <= vector2(0);
	wire_man_prod_w_vector2_range4289w(0) <= vector2(10);
	wire_man_prod_w_vector2_range4299w(0) <= vector2(11);
	wire_man_prod_w_vector2_range4309w(0) <= vector2(12);
	wire_man_prod_w_vector2_range4319w(0) <= vector2(13);
	wire_man_prod_w_vector2_range4329w(0) <= vector2(14);
	wire_man_prod_w_vector2_range4339w(0) <= vector2(15);
	wire_man_prod_w_vector2_range4349w(0) <= vector2(16);
	wire_man_prod_w_vector2_range4359w(0) <= vector2(17);
	wire_man_prod_w_vector2_range4369w(0) <= vector2(18);
	wire_man_prod_w_vector2_range4379w(0) <= vector2(19);
	wire_man_prod_w_vector2_range4199w(0) <= vector2(1);
	wire_man_prod_w_vector2_range4389w(0) <= vector2(20);
	wire_man_prod_w_vector2_range4399w(0) <= vector2(21);
	wire_man_prod_w_vector2_range4409w(0) <= vector2(22);
	wire_man_prod_w_vector2_range4419w(0) <= vector2(23);
	wire_man_prod_w_vector2_range4429w(0) <= vector2(24);
	wire_man_prod_w_vector2_range4439w(0) <= vector2(25);
	wire_man_prod_w_vector2_range4449w(0) <= vector2(26);
	wire_man_prod_w_vector2_range4459w(0) <= vector2(27);
	wire_man_prod_w_vector2_range4469w(0) <= vector2(28);
	wire_man_prod_w_vector2_range4479w(0) <= vector2(29);
	wire_man_prod_w_vector2_range4209w(0) <= vector2(2);
	wire_man_prod_w_vector2_range4489w(0) <= vector2(30);
	wire_man_prod_w_vector2_range4499w(0) <= vector2(31);
	wire_man_prod_w_vector2_range4509w(0) <= vector2(32);
	wire_man_prod_w_vector2_range4519w(0) <= vector2(33);
	wire_man_prod_w_vector2_range4529w(0) <= vector2(34);
	wire_man_prod_w_vector2_range4539w(0) <= vector2(35);
	wire_man_prod_w_vector2_range4549w(0) <= vector2(36);
	wire_man_prod_w_vector2_range4559w(0) <= vector2(37);
	wire_man_prod_w_vector2_range4569w(0) <= vector2(38);
	wire_man_prod_w_vector2_range4579w(0) <= vector2(39);
	wire_man_prod_w_vector2_range4219w(0) <= vector2(3);
	wire_man_prod_w_vector2_range4589w(0) <= vector2(40);
	wire_man_prod_w_vector2_range4599w(0) <= vector2(41);
	wire_man_prod_w_vector2_range4609w(0) <= vector2(42);
	wire_man_prod_w_vector2_range4619w(0) <= vector2(43);
	wire_man_prod_w_vector2_range4629w(0) <= vector2(44);
	wire_man_prod_w_vector2_range4639w(0) <= vector2(45);
	wire_man_prod_w_vector2_range4649w(0) <= vector2(46);
	wire_man_prod_w_vector2_range4659w(0) <= vector2(47);
	wire_man_prod_w_vector2_range4669w(0) <= vector2(48);
	wire_man_prod_w_vector2_range4679w(0) <= vector2(49);
	wire_man_prod_w_vector2_range4229w(0) <= vector2(4);
	wire_man_prod_w_vector2_range4689w(0) <= vector2(50);
	wire_man_prod_w_vector2_range4699w(0) <= vector2(51);
	wire_man_prod_w_vector2_range4709w(0) <= vector2(52);
	wire_man_prod_w_vector2_range4719w(0) <= vector2(53);
	wire_man_prod_w_vector2_range4729w(0) <= vector2(54);
	wire_man_prod_w_vector2_range4739w(0) <= vector2(55);
	wire_man_prod_w_vector2_range4749w(0) <= vector2(56);
	wire_man_prod_w_vector2_range4759w(0) <= vector2(57);
	wire_man_prod_w_vector2_range4769w(0) <= vector2(58);
	wire_man_prod_w_vector2_range4779w(0) <= vector2(59);
	wire_man_prod_w_vector2_range4239w(0) <= vector2(5);
	wire_man_prod_w_vector2_range4789w(0) <= vector2(60);
	wire_man_prod_w_vector2_range4799w(0) <= vector2(61);
	wire_man_prod_w_vector2_range4809w(0) <= vector2(62);
	wire_man_prod_w_vector2_range4819w(0) <= vector2(63);
	wire_man_prod_w_vector2_range4829w(0) <= vector2(64);
	wire_man_prod_w_vector2_range4839w(0) <= vector2(65);
	wire_man_prod_w_vector2_range4849w(0) <= vector2(66);
	wire_man_prod_w_vector2_range4859w(0) <= vector2(67);
	wire_man_prod_w_vector2_range4869w(0) <= vector2(68);
	wire_man_prod_w_vector2_range4879w(0) <= vector2(69);
	wire_man_prod_w_vector2_range4249w(0) <= vector2(6);
	wire_man_prod_w_vector2_range4889w(0) <= vector2(70);
	wire_man_prod_w_vector2_range4899w(0) <= vector2(71);
	wire_man_prod_w_vector2_range4909w(0) <= vector2(72);
	wire_man_prod_w_vector2_range4919w(0) <= vector2(73);
	wire_man_prod_w_vector2_range4929w(0) <= vector2(74);
	wire_man_prod_w_vector2_range4939w(0) <= vector2(75);
	wire_man_prod_w_vector2_range4949w(0) <= vector2(76);
	wire_man_prod_w_vector2_range4959w(0) <= vector2(77);
	wire_man_prod_w_vector2_range4969w(0) <= vector2(78);
	wire_man_prod_w_vector2_range4979w(0) <= vector2(79);
	wire_man_prod_w_vector2_range4259w(0) <= vector2(7);
	wire_man_prod_w_vector2_range4989w(0) <= vector2(80);
	wire_man_prod_w_vector2_range4999w(0) <= vector2(81);
	wire_man_prod_w_vector2_range5009w(0) <= vector2(82);
	wire_man_prod_w_vector2_range5019w(0) <= vector2(83);
	wire_man_prod_w_vector2_range5029w(0) <= vector2(84);
	wire_man_prod_w_vector2_range5039w(0) <= vector2(85);
	wire_man_prod_w_vector2_range5049w(0) <= vector2(86);
	wire_man_prod_w_vector2_range5059w(0) <= vector2(87);
	wire_man_prod_w_vector2_range5069w(0) <= vector2(88);
	wire_man_prod_w_vector2_range5079w(0) <= vector2(89);
	wire_man_prod_w_vector2_range4269w(0) <= vector2(8);
	wire_man_prod_w_vector2_range4279w(0) <= vector2(9);
	sum :  ALTFP_EXa_altmult_opt_csa_ksf
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => car_two_wo,
		datab => sum_two_wo,
		result => wire_sum_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN car_two_adj_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN car_two_adj_reg0 <= car_two_adj;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg0 <= lowest_bits_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg1 <= lowest_bits_wi_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lsb_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lsb_prod_wi_reg0 <= lsb_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mid_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mid_prod_wi_reg0 <= mid_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN msb_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN msb_prod_wi_reg0 <= msb_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sum_two_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sum_two_reg0 <= sum_two;
			END IF;
		END IF;
	END PROCESS;
	compress_a :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 30
	  )
	  PORT MAP ( 
		cout => wire_compress_a_cout,
		dataa => wire_a(59 DOWNTO 30),
		datab => wire_a(29 DOWNTO 0),
		result => wire_compress_a_result
	  );
	compress_b :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 30
	  )
	  PORT MAP ( 
		cout => wire_compress_b_cout,
		dataa => wire_b(59 DOWNTO 30),
		datab => wire_b(29 DOWNTO 0),
		result => wire_compress_b_result
	  );
	lsb_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 30,
		LPM_WIDTHB => 30,
		LPM_WIDTHP => 60,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_a(29 DOWNTO 0),
		datab => wire_b(29 DOWNTO 0),
		result => wire_lsb_prod_result
	  );
	wire_mid_prod_dataa <= ( wire_compress_a_cout & wire_compress_a_result);
	wire_mid_prod_datab <= ( wire_compress_b_cout & wire_compress_b_result);
	mid_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 31,
		LPM_WIDTHB => 31,
		LPM_WIDTHP => 62,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_mid_prod_dataa,
		datab => wire_mid_prod_datab,
		result => wire_mid_prod_result
	  );
	msb_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 30,
		LPM_WIDTHB => 30,
		LPM_WIDTHP => 60,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_a(59 DOWNTO 30),
		datab => wire_b(59 DOWNTO 30),
		result => wire_msb_prod_result
	  );

 END RTL; --ALTFP_EXa_altmult_opt_v4e


--altmult_opt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" LPM_PIPELINE=5 LPM_WIDTHA=61 LPM_WIDTHB=61 LPM_WIDTHP=122 aclr clken clock dataa datab result
--VERSION_BEGIN 16.0 cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END


--altmult_opt_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=2 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=92 aclr clken clock dataa datab result
--VERSION_BEGIN 16.0 cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altmult_opt_csa_nsf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (91 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (91 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (91 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altmult_opt_csa_nsf;

 ARCHITECTURE RTL OF ALTFP_EXa_altmult_opt_csa_nsf IS

	 SIGNAL  wire_add_sub2_result	:	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub2_result;
	add_sub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 92
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub2_result
	  );

 END RTL; --ALTFP_EXa_altmult_opt_csa_nsf

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 lpm_mult 3 reg 464 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altmult_opt_45e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (60 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (60 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (121 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altmult_opt_45e;

 ARCHITECTURE RTL OF ALTFP_EXa_altmult_opt_45e IS

	 SIGNAL  wire_sum_result	:	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL	 car_two_adj_reg0	:	STD_LOGIC_VECTOR(91 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg0	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg1	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg2	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lsb_prod_wi_reg0	:	STD_LOGIC_VECTOR(61 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mid_prod_wi_reg0	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 msb_prod_wi_reg0	:	STD_LOGIC_VECTOR(60 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sum_two_reg0	:	STD_LOGIC_VECTOR(91 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_compress_a_cout	:	STD_LOGIC;
	 SIGNAL  wire_compress_a_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_compress_a_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_compress_b_cout	:	STD_LOGIC;
	 SIGNAL  wire_compress_b_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_compress_b_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_lsb_prod_result	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_mid_prod_dataa	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_mid_prod_datab	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_mid_prod_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_msb_prod_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_msb_prod_result	:	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6615w6624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6555w6725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6549w6735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6543w6745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6537w6755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6531w6765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6525w6775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6519w6785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6513w6795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6507w6805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6501w6815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6609w6635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6495w6825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6489w6835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6483w6845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6477w6855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6471w6865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6465w6875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6459w6885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6453w6895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6447w6905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6441w6915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6603w6645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6435w6925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6429w6935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6423w6945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6417w6955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6411w6965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6405w6975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6399w6985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6393w6995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6387w7005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6381w7015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6597w6655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6375w7025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6369w7035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6363w7045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6357w7055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6351w7065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6345w7075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6339w7085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6333w7095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6327w7105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6321w7115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6591w6665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6315w7125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6309w7135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6303w7145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6297w7155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6291w7165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6285w7175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6279w7185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6273w7195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6267w7205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6261w7215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6585w6675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6255w7225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6248w7235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6244w7245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6240w7255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6236w7265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6232w7275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6228w7285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6224w7295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6220w7305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6216w7315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6579w6685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6212w7325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6208w7335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6204w7345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6200w7355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6196w7365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6192w7375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6188w7385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6184w7395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6180w7405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6176w7415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6573w6695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6172w7425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6168w7435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6164w7445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6160w7455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6156w7465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6152w7475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6148w7485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6144w7495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6140w7505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6136w7515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6567w6705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6132w7525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6126w7535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6561w6715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6622w7551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6724w7662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6734w7673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6744w7684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6754w7695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6764w7706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6774w7717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6784w7728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6794w7739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6804w7750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6814w7761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6634w7563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6824w7772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6834w7783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6844w7794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6854w7805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6864w7816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6874w7827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6884w7838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6894w7849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6904w7860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6914w7871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6644w7574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6924w7882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6934w7893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6944w7904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6954w7915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6964w7926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6974w7937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6984w7948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6994w7959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7004w7970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7014w7981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6654w7585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7024w7992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7034w8003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7044w8014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7054w8025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7064w8036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7074w8047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7084w8058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7094w8069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7104w8080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7114w8091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6664w7596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7124w8102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7134w8113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7144w8124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7154w8135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7164w8146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7174w8157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7184w8168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7194w8179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7204w8190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7214w8201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6674w7607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7224w8212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7234w8223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7244w8234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7254w8245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7264w8256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7274w8267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7284w8278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7294w8289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7304w8300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7314w8311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6684w7618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7324w8322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7334w8333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7344w8344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7354w8355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7364w8366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7374w8377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7384w8388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7394w8399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7404w8410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7414w8421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6694w7629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7424w8432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7434w8443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7444w8454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7454w8465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7464w8476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7474w8487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7484w8498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7494w8509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7504w8520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7514w8531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6704w7640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7524w8542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7534w8553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6714w7651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6616w6617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6556w6557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6550w6551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6544w6545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6538w6539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6532w6533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6526w6527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6520w6521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6514w6515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6508w6509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6502w6503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6610w6611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6496w6497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6490w6491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6484w6485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6478w6479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6472w6473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6466w6467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6460w6461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6454w6455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6448w6449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6442w6443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6604w6605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6436w6437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6430w6431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6424w6425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6418w6419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6412w6413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6406w6407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6400w6401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6394w6395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6388w6389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6382w6383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6598w6599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6376w6377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6370w6371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6364w6365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6358w6359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6352w6353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6346w6347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6340w6341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6334w6335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6328w6329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6322w6323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6592w6593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6316w6317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6310w6311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6304w6305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6298w6299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6292w6293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6286w6287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6280w6281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6274w6275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6268w6269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6262w6263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6586w6587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6256w6257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6250w6251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6580w6581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6574w6575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6568w6569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6562w6563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6613w6614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6553w6554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6547w6548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6541w6542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6535w6536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6529w6530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6523w6524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6517w6518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6511w6512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6505w6506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6499w6500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6607w6608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6493w6494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6487w6488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6481w6482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6475w6476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6469w6470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6463w6464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6457w6458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6451w6452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6445w6446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6439w6440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6601w6602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6433w6434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6427w6428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6421w6422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6415w6416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6409w6410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6403w6404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6397w6398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6391w6392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6385w6386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6379w6380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6595w6596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6373w6374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6367w6368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6361w6362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6355w6356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6349w6350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6343w6344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6337w6338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6331w6332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6325w6326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6319w6320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6589w6590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6313w6314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6307w6308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6301w6302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6295w6296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6289w6290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6283w6284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6277w6278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6271w6272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6265w6266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6259w6260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6583w6584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6253w6254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6577w6578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6571w6572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6565w6566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6559w6560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7546w7553w7554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7658w7664w7665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7669w7675w7676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7680w7686w7687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7691w7697w7698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7702w7708w7709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7713w7719w7720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7724w7730w7731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7735w7741w7742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7746w7752w7753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7757w7763w7764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7559w7565w7566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7768w7774w7775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7779w7785w7786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7790w7796w7797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7801w7807w7808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7812w7818w7819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7823w7829w7830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7834w7840w7841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7845w7851w7852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7856w7862w7863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7867w7873w7874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7570w7576w7577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7878w7884w7885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7889w7895w7896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7900w7906w7907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7911w7917w7918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7922w7928w7929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7933w7939w7940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7944w7950w7951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7955w7961w7962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7966w7972w7973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7977w7983w7984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7581w7587w7588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7988w7994w7995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7999w8005w8006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8010w8016w8017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8021w8027w8028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8032w8038w8039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8043w8049w8050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8054w8060w8061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8065w8071w8072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8076w8082w8083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8087w8093w8094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7592w7598w7599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8098w8104w8105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8109w8115w8116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8120w8126w8127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8131w8137w8138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8142w8148w8149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8153w8159w8160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8164w8170w8171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8175w8181w8182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8186w8192w8193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8197w8203w8204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7603w7609w7610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8208w8214w8215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8219w8225w8226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8230w8236w8237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8241w8247w8248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8252w8258w8259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8263w8269w8270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8274w8280w8281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8285w8291w8292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8296w8302w8303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8307w8313w8314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7614w7620w7621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8318w8324w8325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8329w8335w8336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8340w8346w8347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8351w8357w8358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8362w8368w8369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8373w8379w8380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8384w8390w8391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8395w8401w8402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8406w8412w8413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8417w8423w8424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7625w7631w7632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8428w8434w8435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8439w8445w8446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8450w8456w8457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8461w8467w8468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8472w8478w8479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8483w8489w8490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8494w8500w8501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8505w8511w8512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8516w8522w8523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8527w8533w8534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7636w7642w7643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8538w8544w8545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8549w8555w8556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7647w7653w7654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6619w6626w6627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6721w6727w6728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6731w6737w6738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6741w6747w6748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6751w6757w6758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6761w6767w6768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6771w6777w6778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6781w6787w6788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6791w6797w6798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6801w6807w6808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6811w6817w6818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6631w6637w6638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6821w6827w6828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6831w6837w6838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6841w6847w6848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6851w6857w6858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6861w6867w6868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6871w6877w6878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6881w6887w6888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6891w6897w6898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6901w6907w6908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6911w6917w6918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6641w6647w6648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6921w6927w6928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6931w6937w6938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6941w6947w6948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6951w6957w6958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6961w6967w6968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6971w6977w6978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6981w6987w6988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6991w6997w6998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7001w7007w7008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7011w7017w7018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6651w6657w6658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7021w7027w7028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7031w7037w7038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7041w7047w7048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7051w7057w7058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7061w7067w7068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7071w7077w7078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7081w7087w7088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7091w7097w7098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7101w7107w7108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7111w7117w7118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6661w6667w6668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7121w7127w7128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7131w7137w7138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7141w7147w7148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7151w7157w7158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7161w7167w7168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7171w7177w7178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7181w7187w7188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7191w7197w7198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7201w7207w7208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7211w7217w7218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6671w6677w6678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7221w7227w7228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7231w7237w7238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7241w7247w7248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7251w7257w7258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7261w7267w7268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7271w7277w7278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7281w7287w7288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7291w7297w7298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7301w7307w7308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7311w7317w7318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6681w6687w6688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7321w7327w7328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7331w7337w7338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7341w7347w7348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7351w7357w7358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7361w7367w7368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7371w7377w7378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7381w7387w7388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7391w7397w7398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7401w7407w7408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7411w7417w7418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6691w6697w6698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7421w7427w7428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7431w7437w7438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7441w7447w7448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7451w7457w7458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7461w7467w7468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7471w7477w7478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7481w7487w7488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7491w7497w7498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7501w7507w7508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7511w7517w7518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6701w6707w6708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7521w7527w7528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7531w7537w7538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6711w6717w6718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7546w7553w7554w7555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7658w7664w7665w7666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7669w7675w7676w7677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7680w7686w7687w7688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7691w7697w7698w7699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7702w7708w7709w7710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7713w7719w7720w7721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7724w7730w7731w7732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7735w7741w7742w7743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7746w7752w7753w7754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7757w7763w7764w7765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7559w7565w7566w7567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7768w7774w7775w7776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7779w7785w7786w7787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7790w7796w7797w7798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7801w7807w7808w7809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7812w7818w7819w7820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7823w7829w7830w7831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7834w7840w7841w7842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7845w7851w7852w7853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7856w7862w7863w7864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7867w7873w7874w7875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7570w7576w7577w7578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7878w7884w7885w7886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7889w7895w7896w7897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7900w7906w7907w7908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7911w7917w7918w7919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7922w7928w7929w7930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7933w7939w7940w7941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7944w7950w7951w7952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7955w7961w7962w7963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7966w7972w7973w7974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7977w7983w7984w7985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7581w7587w7588w7589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7988w7994w7995w7996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7999w8005w8006w8007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8010w8016w8017w8018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8021w8027w8028w8029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8032w8038w8039w8040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8043w8049w8050w8051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8054w8060w8061w8062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8065w8071w8072w8073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8076w8082w8083w8084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8087w8093w8094w8095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7592w7598w7599w7600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8098w8104w8105w8106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8109w8115w8116w8117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8120w8126w8127w8128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8131w8137w8138w8139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8142w8148w8149w8150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8153w8159w8160w8161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8164w8170w8171w8172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8175w8181w8182w8183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8186w8192w8193w8194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8197w8203w8204w8205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7603w7609w7610w7611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8208w8214w8215w8216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8219w8225w8226w8227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8230w8236w8237w8238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8241w8247w8248w8249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8252w8258w8259w8260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8263w8269w8270w8271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8274w8280w8281w8282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8285w8291w8292w8293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8296w8302w8303w8304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8307w8313w8314w8315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7614w7620w7621w7622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8318w8324w8325w8326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8329w8335w8336w8337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8340w8346w8347w8348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8351w8357w8358w8359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8362w8368w8369w8370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8373w8379w8380w8381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8384w8390w8391w8392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8395w8401w8402w8403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8406w8412w8413w8414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8417w8423w8424w8425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7625w7631w7632w7633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8428w8434w8435w8436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8439w8445w8446w8447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8450w8456w8457w8458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8461w8467w8468w8469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8472w8478w8479w8480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8483w8489w8490w8491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8494w8500w8501w8502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8505w8511w8512w8513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8516w8522w8523w8524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8527w8533w8534w8535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7636w7642w7643w7644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8538w8544w8545w8546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8549w8555w8556w8557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7647w7653w7654w7655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6619w6626w6627w6628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6721w6727w6728w6729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6731w6737w6738w6739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6741w6747w6748w6749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6751w6757w6758w6759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6761w6767w6768w6769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6771w6777w6778w6779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6781w6787w6788w6789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6791w6797w6798w6799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6801w6807w6808w6809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6811w6817w6818w6819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6631w6637w6638w6639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6821w6827w6828w6829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6831w6837w6838w6839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6841w6847w6848w6849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6851w6857w6858w6859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6861w6867w6868w6869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6871w6877w6878w6879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6881w6887w6888w6889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6891w6897w6898w6899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6901w6907w6908w6909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6911w6917w6918w6919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6641w6647w6648w6649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6921w6927w6928w6929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6931w6937w6938w6939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6941w6947w6948w6949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6951w6957w6958w6959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6961w6967w6968w6969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6971w6977w6978w6979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6981w6987w6988w6989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6991w6997w6998w6999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7001w7007w7008w7009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7011w7017w7018w7019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6651w6657w6658w6659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7021w7027w7028w7029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7031w7037w7038w7039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7041w7047w7048w7049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7051w7057w7058w7059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7061w7067w7068w7069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7071w7077w7078w7079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7081w7087w7088w7089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7091w7097w7098w7099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7101w7107w7108w7109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7111w7117w7118w7119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6661w6667w6668w6669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7121w7127w7128w7129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7131w7137w7138w7139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7141w7147w7148w7149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7151w7157w7158w7159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7161w7167w7168w7169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7171w7177w7178w7179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7181w7187w7188w7189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7191w7197w7198w7199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7201w7207w7208w7209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7211w7217w7218w7219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6671w6677w6678w6679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7221w7227w7228w7229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7231w7237w7238w7239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7241w7247w7248w7249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7251w7257w7258w7259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7261w7267w7268w7269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7271w7277w7278w7279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7281w7287w7288w7289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7291w7297w7298w7299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7301w7307w7308w7309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7311w7317w7318w7319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6681w6687w6688w6689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7321w7327w7328w7329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7331w7337w7338w7339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7341w7347w7348w7349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7351w7357w7358w7359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7361w7367w7368w7369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7371w7377w7378w7379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7381w7387w7388w7389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7391w7397w7398w7399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7401w7407w7408w7409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7411w7417w7418w7419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6691w6697w6698w6699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7421w7427w7428w7429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7431w7437w7438w7439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7441w7447w7448w7449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7451w7457w7458w7459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7461w7467w7468w7469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7471w7477w7478w7479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7481w7487w7488w7489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7491w7497w7498w7499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7501w7507w7508w7509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7511w7517w7518w7519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6701w6707w6708w6709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7521w7527w7528w7529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7531w7537w7538w7539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6711w6717w6718w6719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7546w7547w7548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7658w7659w7660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7669w7670w7671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7680w7681w7682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7691w7692w7693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7702w7703w7704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7713w7714w7715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7724w7725w7726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7735w7736w7737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7746w7747w7748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7757w7758w7759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7559w7560w7561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7768w7769w7770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7779w7780w7781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7790w7791w7792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7801w7802w7803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7812w7813w7814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7823w7824w7825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7834w7835w7836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7845w7846w7847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7856w7857w7858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7867w7868w7869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7570w7571w7572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7878w7879w7880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7889w7890w7891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7900w7901w7902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7911w7912w7913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7922w7923w7924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7933w7934w7935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7944w7945w7946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7955w7956w7957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7966w7967w7968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7977w7978w7979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7581w7582w7583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7988w7989w7990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7999w8000w8001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8010w8011w8012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8021w8022w8023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8032w8033w8034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8043w8044w8045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8054w8055w8056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8065w8066w8067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8076w8077w8078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8087w8088w8089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7592w7593w7594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8098w8099w8100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8109w8110w8111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8120w8121w8122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8131w8132w8133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8142w8143w8144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8153w8154w8155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8164w8165w8166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8175w8176w8177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8186w8187w8188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8197w8198w8199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7603w7604w7605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8208w8209w8210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8219w8220w8221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8230w8231w8232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8241w8242w8243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8252w8253w8254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8263w8264w8265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8274w8275w8276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8285w8286w8287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8296w8297w8298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8307w8308w8309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7614w7615w7616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8318w8319w8320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8329w8330w8331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8340w8341w8342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8351w8352w8353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8362w8363w8364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8373w8374w8375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8384w8385w8386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8395w8396w8397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8406w8407w8408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8417w8418w8419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7625w7626w7627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8428w8429w8430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8439w8440w8441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8450w8451w8452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8461w8462w8463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8472w8473w8474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8483w8484w8485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8494w8495w8496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8505w8506w8507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8516w8517w8518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8527w8528w8529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7636w7637w7638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8538w8539w8540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8549w8550w8551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7647w7648w7649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6619w6620w6621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6721w6722w6723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6731w6732w6733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6741w6742w6743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6751w6752w6753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6761w6762w6763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6771w6772w6773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6781w6782w6783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6791w6792w6793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6801w6802w6803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6811w6812w6813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6631w6632w6633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6821w6822w6823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6831w6832w6833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6841w6842w6843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6851w6852w6853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6861w6862w6863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6871w6872w6873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6881w6882w6883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6891w6892w6893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6901w6902w6903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6911w6912w6913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6641w6642w6643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6921w6922w6923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6931w6932w6933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6941w6942w6943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6951w6952w6953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6961w6962w6963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6971w6972w6973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6981w6982w6983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6991w6992w6993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7001w7002w7003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7011w7012w7013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6651w6652w6653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7021w7022w7023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7031w7032w7033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7041w7042w7043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7051w7052w7053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7061w7062w7063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7071w7072w7073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7081w7082w7083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7091w7092w7093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7101w7102w7103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7111w7112w7113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6661w6662w6663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7121w7122w7123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7131w7132w7133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7141w7142w7143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7151w7152w7153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7161w7162w7163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7171w7172w7173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7181w7182w7183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7191w7192w7193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7201w7202w7203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7211w7212w7213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6671w6672w6673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7221w7222w7223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7231w7232w7233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7241w7242w7243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7251w7252w7253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7261w7262w7263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7271w7272w7273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7281w7282w7283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7291w7292w7293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7301w7302w7303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7311w7312w7313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6681w6682w6683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7321w7322w7323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7331w7332w7333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7341w7342w7343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7351w7352w7353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7361w7362w7363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7371w7372w7373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7381w7382w7383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7391w7392w7393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7401w7402w7403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7411w7412w7413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6691w6692w6693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7421w7422w7423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7431w7432w7433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7441w7442w7443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7451w7452w7453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7461w7462w7463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7471w7472w7473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7481w7482w7483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7491w7492w7493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7501w7502w7503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7511w7512w7513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6701w6702w6703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7521w7522w7523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7531w7532w7533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6711w6712w6713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  car_one :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  car_one_adj :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  car_two :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  car_two_adj :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  car_two_wo :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  lowest_bits_wi :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lowest_bits_wo :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lsb_prod_wi :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  lsb_prod_wo :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  mid_prod_wi :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  mid_prod_wo :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  msb_prod_out :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  msb_prod_wi :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  msb_prod_wo :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  neg_lsb :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  neg_msb :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  sum_one :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  sum_two :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  sum_two_wo :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  vector1 :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  vector2 :	STD_LOGIC_VECTOR (91 DOWNTO 0);
	 SIGNAL  wire_a :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  wire_b :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range8548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_car_one_adj_range7646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_msb_prod_wo_range6559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_lsb_range6564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_neg_msb_range6561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range7534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_sum_one_range6714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range8549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector1_range7647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range7531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_w_vector2_range6711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  ALTFP_EXa_altmult_opt_csa_nsf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(91 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(91 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(91 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6615w6624w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6615w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6618w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6555w6725w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6555w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6558w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6549w6735w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6549w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6552w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6543w6745w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6543w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6546w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6537w6755w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6537w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6540w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6531w6765w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6531w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6534w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6525w6775w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6525w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6528w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6519w6785w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6519w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6522w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6513w6795w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6513w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6516w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6507w6805w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6507w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6510w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6501w6815w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6501w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6609w6635w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6609w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6612w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6495w6825w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6495w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6498w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6489w6835w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6489w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6492w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6483w6845w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6483w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6486w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6477w6855w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6477w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6480w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6471w6865w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6471w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6474w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6465w6875w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6465w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6468w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6459w6885w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6459w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6462w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6453w6895w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6453w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6456w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6447w6905w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6447w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6450w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6441w6915w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6441w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6444w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6603w6645w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6603w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6606w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6435w6925w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6435w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6438w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6429w6935w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6429w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6432w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6423w6945w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6423w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6426w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6417w6955w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6417w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6420w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6411w6965w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6411w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6414w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6405w6975w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6405w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6408w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6399w6985w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6399w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6402w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6393w6995w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6393w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6396w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6387w7005w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6387w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6390w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6381w7015w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6381w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6384w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6597w6655w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6597w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6600w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6375w7025w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6375w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6378w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6369w7035w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6369w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6372w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6363w7045w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6363w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6366w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6357w7055w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6357w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6360w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6351w7065w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6351w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6354w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6345w7075w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6345w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6348w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6339w7085w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6339w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6342w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6333w7095w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6333w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6336w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6327w7105w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6327w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6330w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6321w7115w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6321w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6324w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6591w6665w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6591w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6594w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6315w7125w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6315w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6318w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6309w7135w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6309w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6312w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6303w7145w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6303w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6297w7155w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6297w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6300w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6291w7165w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6291w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6294w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6285w7175w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6285w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6288w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6279w7185w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6279w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6282w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6273w7195w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6273w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6276w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6267w7205w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6267w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6270w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6261w7215w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6261w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6264w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6585w6675w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6585w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6588w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6255w7225w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6255w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6258w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6248w7235w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6248w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6252w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6244w7245w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6244w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6246w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6240w7255w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6240w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6242w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6236w7265w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6236w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6238w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6232w7275w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6232w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6234w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6228w7285w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6228w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6230w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6224w7295w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6224w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6226w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6220w7305w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6220w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6222w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6216w7315w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6216w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6218w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6579w6685w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6579w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6582w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6212w7325w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6212w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6214w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6208w7335w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6208w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6210w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6204w7345w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6204w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6206w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6200w7355w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6200w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6202w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6196w7365w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6196w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6198w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6192w7375w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6192w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6194w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6188w7385w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6188w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6190w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6184w7395w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6184w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6186w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6180w7405w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6180w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6182w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6176w7415w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6176w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6178w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6573w6695w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6573w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6576w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6172w7425w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6172w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6168w7435w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6168w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6170w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6164w7445w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6164w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6166w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6160w7455w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6160w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6162w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6156w7465w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6156w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6158w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6152w7475w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6152w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6154w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6148w7485w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6148w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6150w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6144w7495w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6144w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6146w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6140w7505w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6140w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6142w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6136w7515w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6136w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6138w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6567w6705w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6567w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6570w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6132w7525w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6132w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6134w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6126w7535w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6126w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6129w(0);
	wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6561w6715w(0) <= wire_tbl1_tbl2_prod_w_neg_msb_range6561w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6564w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6622w7551w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6622w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7544w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6724w7662w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6724w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7657w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6734w7673w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6734w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7668w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6744w7684w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6744w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7679w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6754w7695w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6754w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7690w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6764w7706w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6764w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7701w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6774w7717w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6774w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7712w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6784w7728w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6784w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7723w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6794w7739w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6794w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7734w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6804w7750w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6804w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7745w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6814w7761w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6814w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7756w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6634w7563w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6634w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7558w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6824w7772w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6824w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7767w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6834w7783w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6834w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7778w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6844w7794w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6844w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7789w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6854w7805w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6854w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7800w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6864w7816w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6864w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7811w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6874w7827w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6874w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7822w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6884w7838w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6884w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7833w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6894w7849w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6894w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7844w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6904w7860w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6904w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7855w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6914w7871w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6914w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7866w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6644w7574w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6644w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7569w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6924w7882w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6924w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7877w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6934w7893w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6934w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7888w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6944w7904w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6944w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7899w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6954w7915w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6954w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7910w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6964w7926w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6964w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7921w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6974w7937w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6974w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7932w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6984w7948w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6984w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7943w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6994w7959w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6994w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7954w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7004w7970w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7004w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7965w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7014w7981w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7014w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7976w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6654w7585w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6654w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7580w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7024w7992w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7024w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7987w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7034w8003w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7034w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7998w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7044w8014w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7044w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8009w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7054w8025w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7054w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8020w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7064w8036w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7064w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8031w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7074w8047w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7074w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8042w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7084w8058w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7084w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8053w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7094w8069w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7094w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8064w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7104w8080w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7104w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8075w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7114w8091w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7114w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8086w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6664w7596w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6664w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7591w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7124w8102w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7124w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8097w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7134w8113w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7134w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8108w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7144w8124w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7144w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8119w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7154w8135w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7154w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8130w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7164w8146w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7164w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8141w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7174w8157w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7174w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8152w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7184w8168w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7184w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8163w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7194w8179w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7194w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7204w8190w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7204w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8185w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7214w8201w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7214w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8196w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6674w7607w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6674w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7602w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7224w8212w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7224w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8207w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7234w8223w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7234w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8218w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7244w8234w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7244w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8229w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7254w8245w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7254w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8240w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7264w8256w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7264w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8251w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7274w8267w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7274w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8262w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7284w8278w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7284w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8273w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7294w8289w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7294w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8284w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7304w8300w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7304w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8295w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7314w8311w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7314w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6684w7618w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6684w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7613w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7324w8322w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7324w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8317w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7334w8333w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7334w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8328w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7344w8344w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7344w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8339w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7354w8355w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7354w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8350w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7364w8366w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7364w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8361w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7374w8377w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7374w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8372w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7384w8388w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7384w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8383w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7394w8399w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7394w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8394w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7404w8410w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7404w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8405w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7414w8421w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7414w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8416w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6694w7629w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6694w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7624w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7424w8432w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7424w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8427w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7434w8443w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7434w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8438w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7444w8454w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7444w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8449w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7454w8465w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7454w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8460w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7464w8476w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7464w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8471w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7474w8487w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7474w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8482w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7484w8498w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7484w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8493w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7494w8509w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7494w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7504w8520w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7504w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8515w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7514w8531w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7514w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8526w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6704w7640w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6704w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7635w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7524w8542w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7524w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8537w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7534w8553w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range7534w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8548w(0);
	wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6714w7651w(0) <= wire_tbl1_tbl2_prod_w_sum_one_range6714w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7646w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7552w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7546w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7544w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7553w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7546w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6622w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7663w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7658w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7657w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7664w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7658w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6724w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7674w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7669w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7668w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7675w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7669w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6734w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7685w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7680w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7679w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7686w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7680w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6744w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7696w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7691w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7690w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7697w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7691w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6754w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7707w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7702w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7701w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7708w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7702w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6764w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7718w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7713w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7712w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7719w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7713w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6774w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7729w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7724w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7723w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7730w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7724w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6784w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7740w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7735w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7734w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7741w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7735w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6794w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7751w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7746w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7745w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7752w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7746w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6804w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7762w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7757w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7756w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7763w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7757w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6814w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7564w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7559w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7558w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7565w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7559w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6634w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7773w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7768w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7767w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7774w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7768w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6824w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7784w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7779w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7778w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7785w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7779w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6834w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7795w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7790w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7789w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7796w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7790w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6844w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7806w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7801w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7800w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7807w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7801w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6854w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7817w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7812w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7811w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7818w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7812w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6864w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7828w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7823w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7822w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7829w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7823w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6874w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7839w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7834w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7833w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7840w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7834w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6884w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7850w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7845w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7844w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7851w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7845w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6894w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7861w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7856w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7855w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7862w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7856w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6904w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7872w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7867w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7866w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7873w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7867w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6914w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7575w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7570w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7569w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7576w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7570w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6644w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7883w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7878w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7877w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7884w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7878w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6924w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7894w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7889w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7888w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7895w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7889w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6934w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7905w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7900w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7899w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7906w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7900w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6944w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7916w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7911w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7910w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7917w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7911w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6954w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7927w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7922w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7921w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7928w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7922w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6964w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7938w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7933w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7932w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7939w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7933w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6974w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7949w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7944w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7943w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7950w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7944w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6984w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7960w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7955w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7954w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7961w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7955w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6994w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7971w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7966w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7965w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7972w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7966w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7004w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7982w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7977w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7976w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7983w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7977w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7014w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7586w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7581w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7580w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7587w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7581w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6654w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7993w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7988w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7987w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7994w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7988w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7024w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8004w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7999w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7998w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8005w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7999w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7034w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8015w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8010w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8009w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8016w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8010w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7044w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8026w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8021w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8020w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8027w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8021w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7054w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8037w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8032w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8031w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8038w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8032w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7064w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8048w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8043w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8042w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8049w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8043w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7074w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8059w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8054w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8053w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8060w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8054w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7084w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8070w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8065w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8064w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8071w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8065w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7094w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8081w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8076w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8075w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8082w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8076w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7104w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8092w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8087w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8086w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8093w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8087w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7114w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7597w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7592w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7591w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7598w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7592w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6664w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8103w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8098w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8097w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8104w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8098w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7124w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8114w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8109w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8108w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8115w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8109w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7134w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8125w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8120w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8119w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8126w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8120w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7144w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8136w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8131w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8130w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8137w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8131w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7154w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8147w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8142w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8141w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8148w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8142w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7164w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8158w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8153w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8152w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8159w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8153w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8169w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8164w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8163w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8170w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8164w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7184w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8180w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8175w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8181w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8175w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7194w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8191w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8186w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8185w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8192w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8186w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7204w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8202w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8197w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8196w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8203w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8197w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7214w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7608w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7603w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7602w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7609w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7603w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6674w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8213w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8208w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8207w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8214w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8208w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7224w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8224w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8219w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8218w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8225w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8219w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7234w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8235w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8230w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8229w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8236w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8230w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7244w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8246w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8241w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8240w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8247w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8241w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7254w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8257w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8252w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8251w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8258w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8252w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7264w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8268w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8263w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8262w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8269w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8263w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7274w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8279w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8274w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8273w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8280w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8274w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7284w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8290w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8285w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8284w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8291w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8285w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7294w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8301w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8296w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8295w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8302w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8296w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7304w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8312w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8307w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8313w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8307w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7314w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7619w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7614w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7613w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7620w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7614w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6684w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8323w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8318w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8317w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8324w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8318w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7324w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8334w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8329w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8328w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8335w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8329w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7334w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8345w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8340w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8339w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8346w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8340w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7344w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8356w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8351w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8350w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8357w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8351w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7354w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8367w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8362w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8361w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8368w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8362w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7364w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8378w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8373w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8372w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8379w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8373w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7374w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8389w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8384w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8383w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8390w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8384w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7384w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8400w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8395w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8394w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8401w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8395w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7394w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8411w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8406w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8405w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8412w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8406w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7404w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8422w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8417w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8416w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8423w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8417w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7414w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7630w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7625w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7624w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7631w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7625w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6694w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8433w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8428w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8427w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8434w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8428w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7424w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8444w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8439w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8438w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8445w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8439w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7434w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8455w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8450w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8449w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8456w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8450w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7444w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8466w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8461w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8460w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8467w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8461w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7454w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8477w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8472w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8471w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8478w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8472w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7464w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8488w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8483w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8482w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8489w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8483w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7474w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8499w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8494w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8493w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8500w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8494w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7484w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8510w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8505w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8511w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8505w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7494w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8521w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8516w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8515w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8522w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8516w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8532w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8527w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8526w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8533w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8527w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7514w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7641w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7636w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7635w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7642w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7636w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6704w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8543w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8538w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8537w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8544w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8538w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7524w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8554w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8549w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range8548w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8555w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8549w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range7534w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7652w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7647w(0) AND wire_tbl1_tbl2_prod_w_car_one_adj_range7646w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7653w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7647w(0) AND wire_tbl1_tbl2_prod_w_sum_one_range6714w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6625w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6619w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6618w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6626w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6619w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6615w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6726w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6721w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6558w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6727w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6721w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6555w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6736w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6731w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6552w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6737w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6731w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6549w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6746w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6741w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6546w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6747w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6741w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6543w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6756w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6751w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6540w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6757w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6751w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6537w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6766w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6761w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6534w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6767w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6761w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6531w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6776w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6771w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6528w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6777w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6771w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6525w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6786w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6781w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6522w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6787w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6781w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6519w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6796w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6791w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6516w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6797w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6791w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6513w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6806w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6801w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6510w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6807w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6801w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6507w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6816w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6811w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6817w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6811w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6501w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6636w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6631w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6612w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6637w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6631w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6609w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6826w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6821w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6498w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6827w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6821w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6495w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6836w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6831w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6492w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6837w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6831w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6489w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6846w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6841w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6486w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6847w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6841w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6483w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6856w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6851w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6480w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6857w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6851w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6477w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6866w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6861w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6474w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6867w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6861w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6471w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6876w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6871w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6468w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6877w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6871w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6465w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6886w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6881w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6462w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6887w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6881w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6459w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6896w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6891w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6456w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6897w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6891w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6453w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6906w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6901w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6450w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6907w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6901w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6447w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6916w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6911w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6444w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6917w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6911w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6441w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6646w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6641w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6606w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6647w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6641w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6603w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6926w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6921w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6438w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6927w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6921w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6435w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6936w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6931w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6432w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6937w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6931w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6429w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6946w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6941w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6426w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6947w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6941w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6423w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6956w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6951w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6420w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6957w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6951w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6417w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6966w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6961w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6414w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6967w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6961w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6411w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6976w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6971w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6408w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6977w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6971w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6405w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6986w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6981w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6402w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6987w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6981w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6399w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6996w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6991w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6396w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6997w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6991w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6393w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7006w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7001w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6390w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7007w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7001w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6387w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7016w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7011w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6384w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7017w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7011w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6381w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6656w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6651w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6600w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6657w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6651w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6597w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7026w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7021w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6378w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7027w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7021w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6375w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7036w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7031w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6372w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7037w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7031w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6369w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7046w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7041w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6366w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7047w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7041w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6363w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7056w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7051w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6360w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7057w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7051w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6357w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7066w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7061w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6354w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7067w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7061w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6351w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7076w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7071w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6348w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7077w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7071w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6345w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7086w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7081w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6342w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7087w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7081w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6339w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7096w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7091w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6336w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7097w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7091w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6333w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7106w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7101w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6330w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7107w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7101w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6327w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7116w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7111w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6324w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7117w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7111w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6321w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6666w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6661w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6594w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6667w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6661w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6591w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7126w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7121w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6318w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7127w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7121w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6315w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7136w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7131w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6312w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7137w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7131w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6309w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7146w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7141w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7147w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7141w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6303w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7156w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7151w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6300w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7157w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7151w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6297w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7166w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7161w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6294w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7167w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7161w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6291w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7176w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7171w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6288w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7177w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7171w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6285w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7186w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7181w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6282w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7187w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7181w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6279w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7196w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7191w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6276w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7197w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7191w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6273w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7206w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7201w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6270w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7207w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7201w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6267w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7216w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7211w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6264w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7217w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7211w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6261w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6676w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6671w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6588w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6677w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6671w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6585w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7226w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7221w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6258w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7227w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7221w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6255w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7236w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7231w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6252w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7237w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7231w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6248w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7246w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7241w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6246w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7247w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7241w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6244w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7256w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7251w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6242w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7257w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7251w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6240w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7266w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7261w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6238w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7267w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7261w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6236w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7276w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7271w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6234w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7277w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7271w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6232w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7286w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7281w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6230w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7287w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7281w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6228w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7296w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7291w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6226w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7297w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7291w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6224w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7306w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7301w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6222w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7307w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7301w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6220w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7316w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7311w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6218w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7317w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7311w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6216w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6686w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6681w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6582w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6687w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6681w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6579w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7326w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7321w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6214w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7327w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7321w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6212w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7336w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7331w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6210w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7337w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7331w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6208w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7346w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7341w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6206w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7347w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7341w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6204w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7356w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7351w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6202w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7357w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7351w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6200w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7366w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7361w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6198w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7367w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7361w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6196w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7376w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7371w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6194w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7377w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7371w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6192w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7386w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7381w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6190w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7387w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7381w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6188w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7396w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7391w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6186w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7397w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7391w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6184w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7406w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7401w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6182w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7407w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7401w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6180w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7416w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7411w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6178w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7417w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7411w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6176w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6696w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6691w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6576w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6697w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6691w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6573w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7426w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7421w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7427w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7421w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6172w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7436w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7431w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6170w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7437w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7431w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6168w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7446w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7441w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6166w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7447w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7441w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6164w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7456w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7451w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6162w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7457w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7451w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6160w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7466w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7461w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6158w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7467w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7461w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6156w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7476w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7471w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6154w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7477w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7471w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6152w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7486w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7481w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6150w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7487w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7481w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6148w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7496w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7491w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6146w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7497w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7491w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6144w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7506w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7501w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6142w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7507w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7501w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6140w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7516w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7511w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6138w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7517w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7511w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6136w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6706w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6701w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6570w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6707w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6701w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6567w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7526w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7521w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6134w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7527w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7521w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6132w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7536w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7531w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6129w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7537w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7531w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6126w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6716w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6711w(0) AND wire_tbl1_tbl2_prod_w_neg_lsb_range6564w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6717w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6711w(0) AND wire_tbl1_tbl2_prod_w_neg_msb_range6561w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6616w6617w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6616w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6556w6557w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6556w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6550w6551w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6550w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6544w6545w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6544w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6538w6539w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6538w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6532w6533w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6532w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6526w6527w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6526w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6520w6521w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6520w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6514w6515w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6514w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6508w6509w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6508w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6502w6503w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6502w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6610w6611w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6610w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6496w6497w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6496w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6490w6491w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6490w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6484w6485w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6484w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6478w6479w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6478w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6472w6473w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6472w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6466w6467w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6466w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6460w6461w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6460w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6454w6455w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6454w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6448w6449w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6448w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6442w6443w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6442w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6604w6605w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6604w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6436w6437w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6436w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6430w6431w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6430w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6424w6425w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6424w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6418w6419w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6418w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6412w6413w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6412w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6406w6407w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6406w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6400w6401w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6400w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6394w6395w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6394w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6388w6389w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6388w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6382w6383w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6382w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6598w6599w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6598w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6376w6377w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6376w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6370w6371w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6370w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6364w6365w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6364w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6358w6359w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6358w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6352w6353w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6352w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6346w6347w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6346w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6340w6341w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6340w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6334w6335w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6334w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6328w6329w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6328w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6322w6323w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6322w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6592w6593w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6592w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6316w6317w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6316w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6310w6311w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6310w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6304w6305w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6304w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6298w6299w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6298w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6292w6293w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6292w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6286w6287w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6286w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6280w6281w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6280w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6274w6275w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6274w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6268w6269w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6268w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6262w6263w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6262w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6586w6587w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6586w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6256w6257w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6256w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6250w6251w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6250w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6580w6581w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6580w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6574w6575w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6574w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6568w6569w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6568w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6562w6563w(0) <= NOT wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6562w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6613w6614w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6613w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6553w6554w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6553w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6547w6548w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6547w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6541w6542w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6541w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6535w6536w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6535w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6529w6530w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6529w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6523w6524w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6523w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6517w6518w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6517w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6511w6512w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6511w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6505w6506w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6505w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6499w6500w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6499w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6607w6608w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6607w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6493w6494w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6493w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6487w6488w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6487w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6481w6482w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6481w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6475w6476w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6475w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6469w6470w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6469w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6463w6464w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6463w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6457w6458w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6457w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6451w6452w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6451w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6445w6446w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6445w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6439w6440w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6439w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6601w6602w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6601w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6433w6434w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6433w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6427w6428w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6427w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6421w6422w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6421w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6415w6416w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6415w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6409w6410w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6409w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6403w6404w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6403w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6397w6398w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6397w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6391w6392w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6391w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6385w6386w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6385w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6379w6380w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6379w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6595w6596w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6595w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6373w6374w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6373w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6367w6368w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6367w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6361w6362w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6361w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6355w6356w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6355w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6349w6350w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6349w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6343w6344w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6343w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6337w6338w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6337w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6331w6332w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6331w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6325w6326w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6325w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6319w6320w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6319w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6589w6590w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6589w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6313w6314w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6313w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6307w6308w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6307w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6301w6302w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6301w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6295w6296w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6295w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6289w6290w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6289w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6283w6284w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6283w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6277w6278w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6277w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6271w6272w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6271w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6265w6266w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6265w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6259w6260w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6259w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6583w6584w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6583w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6253w6254w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6253w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6577w6578w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6577w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6571w6572w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6571w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6565w6566w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6565w(0);
	wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6559w6560w(0) <= NOT wire_tbl1_tbl2_prod_w_msb_prod_wo_range6559w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7546w7553w7554w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7553w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7552w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7658w7664w7665w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7664w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7663w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7669w7675w7676w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7675w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7674w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7680w7686w7687w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7686w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7685w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7691w7697w7698w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7697w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7696w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7702w7708w7709w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7708w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7707w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7713w7719w7720w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7719w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7718w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7724w7730w7731w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7730w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7729w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7735w7741w7742w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7741w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7740w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7746w7752w7753w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7752w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7751w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7757w7763w7764w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7763w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7762w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7559w7565w7566w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7565w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7564w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7768w7774w7775w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7774w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7773w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7779w7785w7786w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7785w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7784w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7790w7796w7797w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7796w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7795w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7801w7807w7808w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7807w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7806w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7812w7818w7819w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7818w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7817w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7823w7829w7830w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7829w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7828w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7834w7840w7841w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7840w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7839w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7845w7851w7852w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7851w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7850w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7856w7862w7863w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7862w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7861w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7867w7873w7874w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7873w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7872w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7570w7576w7577w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7576w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7575w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7878w7884w7885w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7884w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7883w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7889w7895w7896w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7895w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7894w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7900w7906w7907w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7906w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7905w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7911w7917w7918w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7917w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7916w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7922w7928w7929w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7928w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7927w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7933w7939w7940w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7939w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7938w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7944w7950w7951w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7950w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7949w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7955w7961w7962w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7961w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7960w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7966w7972w7973w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7972w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7971w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7977w7983w7984w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7983w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7982w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7581w7587w7588w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7587w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7586w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7988w7994w7995w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7994w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7993w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7999w8005w8006w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8005w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8004w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8010w8016w8017w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8016w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8015w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8021w8027w8028w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8027w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8026w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8032w8038w8039w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8038w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8037w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8043w8049w8050w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8049w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8048w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8054w8060w8061w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8060w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8059w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8065w8071w8072w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8071w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8070w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8076w8082w8083w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8082w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8081w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8087w8093w8094w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8093w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8092w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7592w7598w7599w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7598w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7597w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8098w8104w8105w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8104w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8103w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8109w8115w8116w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8115w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8114w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8120w8126w8127w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8126w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8125w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8131w8137w8138w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8137w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8136w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8142w8148w8149w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8148w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8147w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8153w8159w8160w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8159w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8158w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8164w8170w8171w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8170w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8169w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8175w8181w8182w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8181w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8180w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8186w8192w8193w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8192w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8191w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8197w8203w8204w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8203w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8202w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7603w7609w7610w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7609w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7608w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8208w8214w8215w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8214w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8213w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8219w8225w8226w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8225w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8224w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8230w8236w8237w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8236w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8235w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8241w8247w8248w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8247w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8246w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8252w8258w8259w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8258w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8257w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8263w8269w8270w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8269w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8268w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8274w8280w8281w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8280w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8279w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8285w8291w8292w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8291w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8290w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8296w8302w8303w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8302w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8301w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8307w8313w8314w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8313w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8312w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7614w7620w7621w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7620w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7619w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8318w8324w8325w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8324w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8323w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8329w8335w8336w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8335w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8334w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8340w8346w8347w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8346w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8345w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8351w8357w8358w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8357w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8356w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8362w8368w8369w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8368w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8367w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8373w8379w8380w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8379w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8378w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8384w8390w8391w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8390w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8389w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8395w8401w8402w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8401w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8400w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8406w8412w8413w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8412w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8411w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8417w8423w8424w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8423w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8422w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7625w7631w7632w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7631w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7630w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8428w8434w8435w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8434w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8433w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8439w8445w8446w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8445w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8444w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8450w8456w8457w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8456w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8455w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8461w8467w8468w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8467w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8466w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8472w8478w8479w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8478w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8477w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8483w8489w8490w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8489w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8488w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8494w8500w8501w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8500w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8499w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8505w8511w8512w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8511w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8510w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8516w8522w8523w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8522w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8521w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8527w8533w8534w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8533w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8532w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7636w7642w7643w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7642w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7641w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8538w8544w8545w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8544w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8543w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8549w8555w8556w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8555w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8554w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7647w7653w7654w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7653w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7652w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6619w6626w6627w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6626w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6625w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6721w6727w6728w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6727w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6726w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6731w6737w6738w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6737w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6736w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6741w6747w6748w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6747w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6746w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6751w6757w6758w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6757w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6756w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6761w6767w6768w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6767w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6766w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6771w6777w6778w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6777w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6776w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6781w6787w6788w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6787w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6786w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6791w6797w6798w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6797w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6796w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6801w6807w6808w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6807w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6806w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6811w6817w6818w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6817w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6816w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6631w6637w6638w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6637w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6636w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6821w6827w6828w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6827w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6826w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6831w6837w6838w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6837w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6836w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6841w6847w6848w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6847w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6846w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6851w6857w6858w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6857w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6856w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6861w6867w6868w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6867w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6866w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6871w6877w6878w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6877w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6876w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6881w6887w6888w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6887w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6886w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6891w6897w6898w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6897w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6896w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6901w6907w6908w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6907w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6906w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6911w6917w6918w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6917w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6916w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6641w6647w6648w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6647w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6646w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6921w6927w6928w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6927w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6926w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6931w6937w6938w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6937w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6936w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6941w6947w6948w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6947w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6946w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6951w6957w6958w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6957w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6956w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6961w6967w6968w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6967w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6966w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6971w6977w6978w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6977w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6976w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6981w6987w6988w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6987w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6986w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6991w6997w6998w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6997w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6996w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7001w7007w7008w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7007w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7006w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7011w7017w7018w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7017w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7016w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6651w6657w6658w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6657w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6656w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7021w7027w7028w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7027w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7026w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7031w7037w7038w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7037w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7036w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7041w7047w7048w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7047w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7046w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7051w7057w7058w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7057w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7056w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7061w7067w7068w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7067w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7066w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7071w7077w7078w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7077w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7076w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7081w7087w7088w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7087w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7086w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7091w7097w7098w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7097w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7096w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7101w7107w7108w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7107w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7106w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7111w7117w7118w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7117w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7116w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6661w6667w6668w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6667w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6666w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7121w7127w7128w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7127w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7126w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7131w7137w7138w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7137w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7136w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7141w7147w7148w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7147w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7146w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7151w7157w7158w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7157w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7156w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7161w7167w7168w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7167w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7166w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7171w7177w7178w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7177w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7176w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7181w7187w7188w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7187w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7186w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7191w7197w7198w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7197w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7196w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7201w7207w7208w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7207w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7206w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7211w7217w7218w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7217w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7216w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6671w6677w6678w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6677w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6676w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7221w7227w7228w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7227w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7226w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7231w7237w7238w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7237w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7236w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7241w7247w7248w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7247w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7246w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7251w7257w7258w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7257w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7256w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7261w7267w7268w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7267w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7266w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7271w7277w7278w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7277w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7276w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7281w7287w7288w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7287w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7286w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7291w7297w7298w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7297w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7296w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7301w7307w7308w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7307w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7311w7317w7318w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7317w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7316w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6681w6687w6688w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6687w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6686w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7321w7327w7328w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7327w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7326w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7331w7337w7338w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7337w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7336w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7341w7347w7348w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7347w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7346w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7351w7357w7358w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7357w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7356w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7361w7367w7368w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7367w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7366w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7371w7377w7378w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7377w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7376w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7381w7387w7388w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7387w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7386w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7391w7397w7398w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7397w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7396w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7401w7407w7408w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7407w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7406w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7411w7417w7418w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7417w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7416w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6691w6697w6698w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6697w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6696w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7421w7427w7428w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7427w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7426w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7431w7437w7438w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7437w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7436w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7441w7447w7448w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7447w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7446w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7451w7457w7458w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7457w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7456w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7461w7467w7468w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7467w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7466w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7471w7477w7478w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7477w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7476w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7481w7487w7488w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7487w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7486w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7491w7497w7498w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7497w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7496w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7501w7507w7508w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7507w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7506w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7511w7517w7518w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7517w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7516w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6701w6707w6708w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6707w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6706w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7521w7527w7528w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7527w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7526w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7531w7537w7538w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7537w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7536w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6711w6717w6718w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6717w(0) OR wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6716w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7546w7553w7554w7555w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7546w7553w7554w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6622w7551w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7658w7664w7665w7666w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7658w7664w7665w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6724w7662w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7669w7675w7676w7677w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7669w7675w7676w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6734w7673w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7680w7686w7687w7688w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7680w7686w7687w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6744w7684w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7691w7697w7698w7699w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7691w7697w7698w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6754w7695w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7702w7708w7709w7710w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7702w7708w7709w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6764w7706w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7713w7719w7720w7721w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7713w7719w7720w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6774w7717w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7724w7730w7731w7732w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7724w7730w7731w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6784w7728w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7735w7741w7742w7743w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7735w7741w7742w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6794w7739w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7746w7752w7753w7754w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7746w7752w7753w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6804w7750w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7757w7763w7764w7765w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7757w7763w7764w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6814w7761w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7559w7565w7566w7567w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7559w7565w7566w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6634w7563w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7768w7774w7775w7776w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7768w7774w7775w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6824w7772w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7779w7785w7786w7787w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7779w7785w7786w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6834w7783w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7790w7796w7797w7798w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7790w7796w7797w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6844w7794w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7801w7807w7808w7809w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7801w7807w7808w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6854w7805w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7812w7818w7819w7820w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7812w7818w7819w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6864w7816w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7823w7829w7830w7831w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7823w7829w7830w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6874w7827w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7834w7840w7841w7842w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7834w7840w7841w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6884w7838w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7845w7851w7852w7853w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7845w7851w7852w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6894w7849w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7856w7862w7863w7864w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7856w7862w7863w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6904w7860w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7867w7873w7874w7875w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7867w7873w7874w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6914w7871w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7570w7576w7577w7578w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7570w7576w7577w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6644w7574w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7878w7884w7885w7886w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7878w7884w7885w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6924w7882w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7889w7895w7896w7897w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7889w7895w7896w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6934w7893w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7900w7906w7907w7908w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7900w7906w7907w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6944w7904w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7911w7917w7918w7919w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7911w7917w7918w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6954w7915w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7922w7928w7929w7930w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7922w7928w7929w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6964w7926w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7933w7939w7940w7941w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7933w7939w7940w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6974w7937w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7944w7950w7951w7952w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7944w7950w7951w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6984w7948w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7955w7961w7962w7963w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7955w7961w7962w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6994w7959w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7966w7972w7973w7974w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7966w7972w7973w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7004w7970w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7977w7983w7984w7985w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7977w7983w7984w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7014w7981w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7581w7587w7588w7589w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7581w7587w7588w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6654w7585w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7988w7994w7995w7996w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7988w7994w7995w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7024w7992w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7999w8005w8006w8007w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7999w8005w8006w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7034w8003w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8010w8016w8017w8018w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8010w8016w8017w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7044w8014w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8021w8027w8028w8029w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8021w8027w8028w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7054w8025w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8032w8038w8039w8040w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8032w8038w8039w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7064w8036w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8043w8049w8050w8051w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8043w8049w8050w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7074w8047w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8054w8060w8061w8062w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8054w8060w8061w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7084w8058w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8065w8071w8072w8073w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8065w8071w8072w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7094w8069w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8076w8082w8083w8084w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8076w8082w8083w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7104w8080w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8087w8093w8094w8095w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8087w8093w8094w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7114w8091w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7592w7598w7599w7600w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7592w7598w7599w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6664w7596w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8098w8104w8105w8106w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8098w8104w8105w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7124w8102w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8109w8115w8116w8117w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8109w8115w8116w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7134w8113w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8120w8126w8127w8128w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8120w8126w8127w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7144w8124w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8131w8137w8138w8139w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8131w8137w8138w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7154w8135w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8142w8148w8149w8150w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8142w8148w8149w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7164w8146w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8153w8159w8160w8161w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8153w8159w8160w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7174w8157w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8164w8170w8171w8172w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8164w8170w8171w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7184w8168w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8175w8181w8182w8183w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8175w8181w8182w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7194w8179w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8186w8192w8193w8194w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8186w8192w8193w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7204w8190w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8197w8203w8204w8205w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8197w8203w8204w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7214w8201w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7603w7609w7610w7611w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7603w7609w7610w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6674w7607w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8208w8214w8215w8216w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8208w8214w8215w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7224w8212w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8219w8225w8226w8227w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8219w8225w8226w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7234w8223w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8230w8236w8237w8238w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8230w8236w8237w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7244w8234w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8241w8247w8248w8249w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8241w8247w8248w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7254w8245w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8252w8258w8259w8260w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8252w8258w8259w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7264w8256w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8263w8269w8270w8271w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8263w8269w8270w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7274w8267w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8274w8280w8281w8282w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8274w8280w8281w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7284w8278w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8285w8291w8292w8293w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8285w8291w8292w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7294w8289w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8296w8302w8303w8304w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8296w8302w8303w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7304w8300w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8307w8313w8314w8315w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8307w8313w8314w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7314w8311w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7614w7620w7621w7622w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7614w7620w7621w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6684w7618w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8318w8324w8325w8326w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8318w8324w8325w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7324w8322w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8329w8335w8336w8337w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8329w8335w8336w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7334w8333w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8340w8346w8347w8348w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8340w8346w8347w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7344w8344w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8351w8357w8358w8359w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8351w8357w8358w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7354w8355w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8362w8368w8369w8370w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8362w8368w8369w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7364w8366w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8373w8379w8380w8381w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8373w8379w8380w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7374w8377w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8384w8390w8391w8392w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8384w8390w8391w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7384w8388w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8395w8401w8402w8403w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8395w8401w8402w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7394w8399w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8406w8412w8413w8414w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8406w8412w8413w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7404w8410w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8417w8423w8424w8425w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8417w8423w8424w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7414w8421w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7625w7631w7632w7633w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7625w7631w7632w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6694w7629w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8428w8434w8435w8436w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8428w8434w8435w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7424w8432w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8439w8445w8446w8447w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8439w8445w8446w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7434w8443w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8450w8456w8457w8458w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8450w8456w8457w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7444w8454w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8461w8467w8468w8469w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8461w8467w8468w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7454w8465w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8472w8478w8479w8480w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8472w8478w8479w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7464w8476w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8483w8489w8490w8491w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8483w8489w8490w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7474w8487w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8494w8500w8501w8502w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8494w8500w8501w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7484w8498w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8505w8511w8512w8513w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8505w8511w8512w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7494w8509w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8516w8522w8523w8524w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8516w8522w8523w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7504w8520w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8527w8533w8534w8535w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8527w8533w8534w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7514w8531w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7636w7642w7643w7644w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7636w7642w7643w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6704w7640w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8538w8544w8545w8546w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8538w8544w8545w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7524w8542w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8549w8555w8556w8557w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8549w8555w8556w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range7534w8553w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7647w7653w7654w7655w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7647w7653w7654w(0) OR wire_tbl1_tbl2_prod_w_lg_w_sum_one_range6714w7651w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6619w6626w6627w6628w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6619w6626w6627w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6615w6624w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6721w6727w6728w6729w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6721w6727w6728w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6555w6725w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6731w6737w6738w6739w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6731w6737w6738w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6549w6735w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6741w6747w6748w6749w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6741w6747w6748w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6543w6745w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6751w6757w6758w6759w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6751w6757w6758w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6537w6755w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6761w6767w6768w6769w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6761w6767w6768w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6531w6765w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6771w6777w6778w6779w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6771w6777w6778w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6525w6775w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6781w6787w6788w6789w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6781w6787w6788w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6519w6785w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6791w6797w6798w6799w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6791w6797w6798w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6513w6795w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6801w6807w6808w6809w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6801w6807w6808w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6507w6805w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6811w6817w6818w6819w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6811w6817w6818w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6501w6815w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6631w6637w6638w6639w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6631w6637w6638w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6609w6635w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6821w6827w6828w6829w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6821w6827w6828w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6495w6825w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6831w6837w6838w6839w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6831w6837w6838w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6489w6835w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6841w6847w6848w6849w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6841w6847w6848w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6483w6845w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6851w6857w6858w6859w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6851w6857w6858w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6477w6855w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6861w6867w6868w6869w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6861w6867w6868w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6471w6865w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6871w6877w6878w6879w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6871w6877w6878w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6465w6875w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6881w6887w6888w6889w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6881w6887w6888w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6459w6885w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6891w6897w6898w6899w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6891w6897w6898w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6453w6895w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6901w6907w6908w6909w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6901w6907w6908w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6447w6905w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6911w6917w6918w6919w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6911w6917w6918w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6441w6915w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6641w6647w6648w6649w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6641w6647w6648w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6603w6645w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6921w6927w6928w6929w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6921w6927w6928w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6435w6925w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6931w6937w6938w6939w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6931w6937w6938w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6429w6935w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6941w6947w6948w6949w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6941w6947w6948w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6423w6945w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6951w6957w6958w6959w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6951w6957w6958w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6417w6955w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6961w6967w6968w6969w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6961w6967w6968w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6411w6965w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6971w6977w6978w6979w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6971w6977w6978w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6405w6975w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6981w6987w6988w6989w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6981w6987w6988w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6399w6985w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6991w6997w6998w6999w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6991w6997w6998w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6393w6995w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7001w7007w7008w7009w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7001w7007w7008w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6387w7005w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7011w7017w7018w7019w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7011w7017w7018w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6381w7015w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6651w6657w6658w6659w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6651w6657w6658w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6597w6655w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7021w7027w7028w7029w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7021w7027w7028w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6375w7025w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7031w7037w7038w7039w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7031w7037w7038w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6369w7035w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7041w7047w7048w7049w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7041w7047w7048w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6363w7045w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7051w7057w7058w7059w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7051w7057w7058w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6357w7055w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7061w7067w7068w7069w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7061w7067w7068w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6351w7065w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7071w7077w7078w7079w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7071w7077w7078w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6345w7075w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7081w7087w7088w7089w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7081w7087w7088w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6339w7085w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7091w7097w7098w7099w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7091w7097w7098w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6333w7095w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7101w7107w7108w7109w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7101w7107w7108w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6327w7105w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7111w7117w7118w7119w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7111w7117w7118w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6321w7115w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6661w6667w6668w6669w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6661w6667w6668w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6591w6665w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7121w7127w7128w7129w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7121w7127w7128w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6315w7125w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7131w7137w7138w7139w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7131w7137w7138w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6309w7135w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7141w7147w7148w7149w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7141w7147w7148w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6303w7145w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7151w7157w7158w7159w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7151w7157w7158w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6297w7155w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7161w7167w7168w7169w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7161w7167w7168w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6291w7165w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7171w7177w7178w7179w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7171w7177w7178w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6285w7175w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7181w7187w7188w7189w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7181w7187w7188w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6279w7185w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7191w7197w7198w7199w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7191w7197w7198w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6273w7195w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7201w7207w7208w7209w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7201w7207w7208w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6267w7205w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7211w7217w7218w7219w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7211w7217w7218w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6261w7215w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6671w6677w6678w6679w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6671w6677w6678w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6585w6675w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7221w7227w7228w7229w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7221w7227w7228w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6255w7225w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7231w7237w7238w7239w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7231w7237w7238w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6248w7235w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7241w7247w7248w7249w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7241w7247w7248w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6244w7245w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7251w7257w7258w7259w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7251w7257w7258w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6240w7255w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7261w7267w7268w7269w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7261w7267w7268w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6236w7265w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7271w7277w7278w7279w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7271w7277w7278w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6232w7275w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7281w7287w7288w7289w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7281w7287w7288w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6228w7285w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7291w7297w7298w7299w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7291w7297w7298w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6224w7295w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7301w7307w7308w7309w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7301w7307w7308w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6220w7305w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7311w7317w7318w7319w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7311w7317w7318w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6216w7315w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6681w6687w6688w6689w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6681w6687w6688w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6579w6685w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7321w7327w7328w7329w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7321w7327w7328w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6212w7325w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7331w7337w7338w7339w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7331w7337w7338w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6208w7335w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7341w7347w7348w7349w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7341w7347w7348w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6204w7345w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7351w7357w7358w7359w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7351w7357w7358w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6200w7355w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7361w7367w7368w7369w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7361w7367w7368w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6196w7365w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7371w7377w7378w7379w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7371w7377w7378w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6192w7375w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7381w7387w7388w7389w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7381w7387w7388w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6188w7385w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7391w7397w7398w7399w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7391w7397w7398w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6184w7395w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7401w7407w7408w7409w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7401w7407w7408w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6180w7405w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7411w7417w7418w7419w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7411w7417w7418w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6176w7415w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6691w6697w6698w6699w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6691w6697w6698w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6573w6695w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7421w7427w7428w7429w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7421w7427w7428w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6172w7425w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7431w7437w7438w7439w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7431w7437w7438w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6168w7435w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7441w7447w7448w7449w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7441w7447w7448w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6164w7445w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7451w7457w7458w7459w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7451w7457w7458w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6160w7455w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7461w7467w7468w7469w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7461w7467w7468w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6156w7465w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7471w7477w7478w7479w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7471w7477w7478w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6152w7475w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7481w7487w7488w7489w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7481w7487w7488w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6148w7485w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7491w7497w7498w7499w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7491w7497w7498w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6144w7495w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7501w7507w7508w7509w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7501w7507w7508w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6140w7505w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7511w7517w7518w7519w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7511w7517w7518w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6136w7515w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6701w6707w6708w6709w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6701w6707w6708w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6567w6705w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7521w7527w7528w7529w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7521w7527w7528w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6132w7525w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7531w7537w7538w7539w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7531w7537w7538w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6126w7535w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6711w6717w6718w6719w(0) <= wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6711w6717w6718w(0) OR wire_tbl1_tbl2_prod_w_lg_w_neg_msb_range6561w6715w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7546w7547w7548w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7547w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7544w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7658w7659w7660w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7659w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7657w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7669w7670w7671w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7670w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7668w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7680w7681w7682w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7681w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7679w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7691w7692w7693w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7692w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7690w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7702w7703w7704w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7703w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7701w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7713w7714w7715w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7714w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7712w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7724w7725w7726w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7725w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7723w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7735w7736w7737w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7736w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7734w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7746w7747w7748w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7747w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7745w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7757w7758w7759w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7758w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7756w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7559w7560w7561w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7560w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7558w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7768w7769w7770w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7769w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7767w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7779w7780w7781w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7780w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7778w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7790w7791w7792w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7791w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7789w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7801w7802w7803w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7802w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7800w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7812w7813w7814w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7813w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7811w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7823w7824w7825w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7824w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7822w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7834w7835w7836w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7835w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7833w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7845w7846w7847w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7846w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7844w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7856w7857w7858w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7857w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7855w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7867w7868w7869w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7868w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7866w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7570w7571w7572w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7571w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7569w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7878w7879w7880w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7879w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7877w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7889w7890w7891w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7890w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7888w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7900w7901w7902w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7901w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7899w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7911w7912w7913w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7912w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7910w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7922w7923w7924w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7923w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7921w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7933w7934w7935w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7934w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7932w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7944w7945w7946w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7945w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7943w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7955w7956w7957w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7956w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7954w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7966w7967w7968w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7967w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7965w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7977w7978w7979w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7978w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7976w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7581w7582w7583w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7582w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7580w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7988w7989w7990w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7989w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7987w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7999w8000w8001w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8000w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7998w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8010w8011w8012w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8011w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8009w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8021w8022w8023w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8022w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8020w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8032w8033w8034w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8033w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8031w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8043w8044w8045w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8044w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8042w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8054w8055w8056w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8055w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8053w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8065w8066w8067w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8066w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8064w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8076w8077w8078w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8077w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8075w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8087w8088w8089w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8088w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8086w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7592w7593w7594w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7593w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7591w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8098w8099w8100w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8099w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8097w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8109w8110w8111w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8110w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8108w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8120w8121w8122w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8121w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8119w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8131w8132w8133w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8132w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8130w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8142w8143w8144w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8143w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8141w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8153w8154w8155w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8154w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8152w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8164w8165w8166w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8165w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8163w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8175w8176w8177w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8176w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8186w8187w8188w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8187w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8185w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8197w8198w8199w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8198w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8196w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7603w7604w7605w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7604w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7602w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8208w8209w8210w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8209w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8207w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8219w8220w8221w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8220w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8218w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8230w8231w8232w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8231w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8229w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8241w8242w8243w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8242w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8240w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8252w8253w8254w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8253w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8251w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8263w8264w8265w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8264w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8262w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8274w8275w8276w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8275w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8273w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8285w8286w8287w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8286w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8284w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8296w8297w8298w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8297w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8295w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8307w8308w8309w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8308w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7614w7615w7616w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7615w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7613w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8318w8319w8320w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8319w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8317w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8329w8330w8331w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8330w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8328w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8340w8341w8342w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8341w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8339w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8351w8352w8353w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8352w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8350w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8362w8363w8364w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8363w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8361w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8373w8374w8375w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8374w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8372w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8384w8385w8386w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8385w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8383w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8395w8396w8397w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8396w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8394w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8406w8407w8408w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8407w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8405w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8417w8418w8419w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8418w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8416w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7625w7626w7627w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7626w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7624w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8428w8429w8430w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8429w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8427w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8439w8440w8441w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8440w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8438w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8450w8451w8452w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8451w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8449w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8461w8462w8463w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8462w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8460w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8472w8473w8474w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8473w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8471w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8483w8484w8485w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8484w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8482w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8494w8495w8496w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8495w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8493w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8505w8506w8507w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8506w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8516w8517w8518w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8517w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8515w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8527w8528w8529w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8528w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8526w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7636w7637w7638w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7637w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7635w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8538w8539w8540w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8539w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8537w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8549w8550w8551w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8550w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range8548w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7647w7648w7649w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7648w(0) XOR wire_tbl1_tbl2_prod_w_car_one_adj_range7646w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6619w6620w6621w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6620w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6618w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6721w6722w6723w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6722w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6558w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6731w6732w6733w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6732w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6552w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6741w6742w6743w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6742w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6546w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6751w6752w6753w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6752w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6540w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6761w6762w6763w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6762w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6534w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6771w6772w6773w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6772w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6528w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6781w6782w6783w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6782w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6522w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6791w6792w6793w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6792w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6516w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6801w6802w6803w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6802w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6510w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6811w6812w6813w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6812w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6631w6632w6633w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6632w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6612w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6821w6822w6823w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6822w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6498w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6831w6832w6833w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6832w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6492w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6841w6842w6843w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6842w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6486w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6851w6852w6853w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6852w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6480w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6861w6862w6863w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6862w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6474w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6871w6872w6873w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6872w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6468w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6881w6882w6883w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6882w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6462w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6891w6892w6893w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6892w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6456w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6901w6902w6903w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6902w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6450w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6911w6912w6913w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6912w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6444w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6641w6642w6643w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6642w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6606w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6921w6922w6923w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6922w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6438w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6931w6932w6933w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6932w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6432w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6941w6942w6943w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6942w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6426w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6951w6952w6953w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6952w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6420w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6961w6962w6963w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6962w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6414w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6971w6972w6973w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6972w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6408w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6981w6982w6983w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6982w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6402w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6991w6992w6993w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6992w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6396w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7001w7002w7003w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7002w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6390w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7011w7012w7013w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7012w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6384w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6651w6652w6653w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6652w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6600w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7021w7022w7023w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7022w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6378w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7031w7032w7033w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7032w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6372w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7041w7042w7043w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7042w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6366w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7051w7052w7053w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7052w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6360w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7061w7062w7063w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7062w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6354w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7071w7072w7073w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7072w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6348w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7081w7082w7083w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7082w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6342w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7091w7092w7093w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7092w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6336w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7101w7102w7103w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7102w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6330w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7111w7112w7113w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7112w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6324w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6661w6662w6663w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6662w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6594w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7121w7122w7123w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7122w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6318w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7131w7132w7133w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7132w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6312w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7141w7142w7143w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7142w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6306w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7151w7152w7153w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7152w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6300w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7161w7162w7163w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7162w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6294w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7171w7172w7173w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7172w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6288w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7181w7182w7183w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7182w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6282w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7191w7192w7193w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7192w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6276w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7201w7202w7203w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7202w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6270w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7211w7212w7213w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7212w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6264w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6671w6672w6673w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6672w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6588w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7221w7222w7223w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7222w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6258w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7231w7232w7233w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7232w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6252w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7241w7242w7243w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7242w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6246w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7251w7252w7253w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7252w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6242w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7261w7262w7263w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7262w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6238w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7271w7272w7273w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7272w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6234w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7281w7282w7283w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7282w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6230w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7291w7292w7293w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7292w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6226w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7301w7302w7303w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7302w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6222w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7311w7312w7313w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7312w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6218w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6681w6682w6683w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6682w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6582w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7321w7322w7323w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7322w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6214w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7331w7332w7333w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7332w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6210w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7341w7342w7343w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7342w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6206w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7351w7352w7353w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7352w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6202w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7361w7362w7363w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7362w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6198w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7371w7372w7373w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7372w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6194w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7381w7382w7383w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7382w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6190w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7391w7392w7393w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7392w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6186w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7401w7402w7403w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7402w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6182w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7411w7412w7413w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7412w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6178w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6691w6692w6693w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6692w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6576w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7421w7422w7423w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7422w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7431w7432w7433w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7432w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6170w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7441w7442w7443w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7442w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6166w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7451w7452w7453w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7452w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6162w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7461w7462w7463w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7462w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6158w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7471w7472w7473w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7472w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6154w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7481w7482w7483w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7482w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6150w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7491w7492w7493w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7492w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6146w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7501w7502w7503w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7502w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6142w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7511w7512w7513w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7512w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6138w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6701w6702w6703w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6702w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6570w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7521w7522w7523w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7522w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6134w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7531w7532w7533w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7532w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6129w(0);
	wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6711w6712w6713w(0) <= wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6712w(0) XOR wire_tbl1_tbl2_prod_w_neg_lsb_range6564w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7546w7547w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7546w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6622w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7658w7659w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7658w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6724w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7669w7670w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7669w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6734w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7680w7681w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7680w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6744w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7691w7692w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7691w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6754w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7702w7703w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7702w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6764w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7713w7714w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7713w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6774w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7724w7725w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7724w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6784w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7735w7736w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7735w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6794w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7746w7747w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7746w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6804w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7757w7758w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7757w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6814w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7559w7560w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7559w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6634w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7768w7769w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7768w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6824w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7779w7780w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7779w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6834w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7790w7791w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7790w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6844w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7801w7802w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7801w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6854w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7812w7813w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7812w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6864w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7823w7824w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7823w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6874w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7834w7835w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7834w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6884w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7845w7846w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7845w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6894w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7856w7857w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7856w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6904w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7867w7868w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7867w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6914w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7570w7571w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7570w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6644w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7878w7879w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7878w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6924w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7889w7890w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7889w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6934w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7900w7901w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7900w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6944w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7911w7912w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7911w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6954w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7922w7923w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7922w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6964w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7933w7934w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7933w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6974w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7944w7945w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7944w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6984w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7955w7956w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7955w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6994w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7966w7967w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7966w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7004w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7977w7978w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7977w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7014w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7581w7582w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7581w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6654w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7988w7989w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7988w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7024w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7999w8000w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7999w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7034w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8010w8011w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8010w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7044w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8021w8022w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8021w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7054w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8032w8033w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8032w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7064w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8043w8044w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8043w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7074w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8054w8055w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8054w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7084w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8065w8066w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8065w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7094w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8076w8077w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8076w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7104w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8087w8088w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8087w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7114w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7592w7593w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7592w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6664w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8098w8099w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8098w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7124w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8109w8110w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8109w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7134w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8120w8121w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8120w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7144w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8131w8132w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8131w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7154w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8142w8143w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8142w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7164w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8153w8154w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8153w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7174w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8164w8165w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8164w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7184w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8175w8176w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8175w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7194w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8186w8187w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8186w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7204w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8197w8198w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8197w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7214w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7603w7604w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7603w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6674w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8208w8209w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8208w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7224w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8219w8220w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8219w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7234w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8230w8231w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8230w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7244w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8241w8242w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8241w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7254w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8252w8253w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8252w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7264w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8263w8264w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8263w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7274w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8274w8275w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8274w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7284w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8285w8286w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8285w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7294w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8296w8297w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8296w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7304w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8307w8308w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8307w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7314w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7614w7615w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7614w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6684w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8318w8319w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8318w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7324w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8329w8330w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8329w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7334w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8340w8341w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8340w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7344w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8351w8352w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8351w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7354w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8362w8363w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8362w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7364w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8373w8374w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8373w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7374w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8384w8385w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8384w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7384w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8395w8396w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8395w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7394w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8406w8407w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8406w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7404w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8417w8418w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8417w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7414w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7625w7626w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7625w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6694w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8428w8429w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8428w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7424w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8439w8440w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8439w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7434w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8450w8451w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8450w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7444w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8461w8462w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8461w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7454w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8472w8473w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8472w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7464w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8483w8484w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8483w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7474w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8494w8495w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8494w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7484w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8505w8506w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8505w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7494w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8516w8517w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8516w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7504w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8527w8528w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8527w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7514w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7636w7637w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7636w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6704w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8538w8539w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8538w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7524w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range8549w8550w(0) <= wire_tbl1_tbl2_prod_w_vector1_range8549w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range7534w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector1_range7647w7648w(0) <= wire_tbl1_tbl2_prod_w_vector1_range7647w(0) XOR wire_tbl1_tbl2_prod_w_sum_one_range6714w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6619w6620w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6619w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6615w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6721w6722w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6721w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6555w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6731w6732w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6731w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6549w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6741w6742w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6741w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6543w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6751w6752w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6751w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6537w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6761w6762w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6761w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6531w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6771w6772w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6771w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6525w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6781w6782w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6781w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6519w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6791w6792w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6791w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6513w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6801w6802w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6801w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6507w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6811w6812w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6811w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6501w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6631w6632w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6631w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6609w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6821w6822w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6821w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6495w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6831w6832w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6831w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6489w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6841w6842w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6841w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6483w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6851w6852w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6851w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6477w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6861w6862w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6861w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6471w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6871w6872w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6871w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6465w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6881w6882w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6881w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6459w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6891w6892w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6891w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6453w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6901w6902w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6901w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6447w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6911w6912w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6911w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6441w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6641w6642w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6641w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6603w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6921w6922w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6921w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6435w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6931w6932w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6931w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6429w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6941w6942w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6941w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6423w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6951w6952w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6951w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6417w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6961w6962w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6961w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6411w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6971w6972w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6971w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6405w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6981w6982w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6981w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6399w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6991w6992w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6991w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6393w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7001w7002w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7001w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6387w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7011w7012w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7011w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6381w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6651w6652w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6651w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6597w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7021w7022w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7021w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6375w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7031w7032w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7031w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6369w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7041w7042w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7041w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6363w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7051w7052w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7051w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6357w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7061w7062w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7061w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6351w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7071w7072w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7071w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6345w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7081w7082w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7081w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6339w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7091w7092w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7091w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6333w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7101w7102w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7101w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6327w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7111w7112w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7111w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6321w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6661w6662w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6661w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6591w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7121w7122w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7121w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6315w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7131w7132w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7131w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6309w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7141w7142w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7141w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6303w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7151w7152w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7151w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6297w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7161w7162w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7161w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6291w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7171w7172w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7171w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6285w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7181w7182w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7181w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6279w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7191w7192w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7191w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6273w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7201w7202w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7201w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6267w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7211w7212w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7211w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6261w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6671w6672w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6671w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6585w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7221w7222w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7221w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6255w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7231w7232w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7231w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6248w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7241w7242w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7241w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6244w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7251w7252w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7251w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6240w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7261w7262w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7261w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6236w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7271w7272w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7271w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6232w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7281w7282w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7281w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6228w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7291w7292w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7291w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6224w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7301w7302w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7301w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6220w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7311w7312w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7311w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6216w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6681w6682w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6681w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6579w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7321w7322w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7321w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6212w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7331w7332w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7331w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6208w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7341w7342w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7341w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6204w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7351w7352w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7351w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6200w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7361w7362w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7361w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6196w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7371w7372w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7371w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6192w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7381w7382w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7381w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6188w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7391w7392w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7391w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6184w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7401w7402w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7401w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6180w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7411w7412w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7411w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6176w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6691w6692w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6691w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6573w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7421w7422w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7421w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6172w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7431w7432w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7431w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6168w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7441w7442w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7441w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6164w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7451w7452w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7451w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6160w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7461w7462w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7461w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6156w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7471w7472w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7471w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6152w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7481w7482w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7481w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6148w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7491w7492w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7491w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6144w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7501w7502w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7501w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6140w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7511w7512w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7511w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6136w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6701w6702w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6701w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6567w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7521w7522w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7521w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6132w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range7531w7532w(0) <= wire_tbl1_tbl2_prod_w_vector2_range7531w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6126w(0);
	wire_tbl1_tbl2_prod_w_lg_w_vector2_range6711w6712w(0) <= wire_tbl1_tbl2_prod_w_vector2_range6711w(0) XOR wire_tbl1_tbl2_prod_w_neg_msb_range6561w(0);
	car_one <= ( wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7531w7537w7538w7539w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7521w7527w7528w7529w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7511w7517w7518w7519w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7501w7507w7508w7509w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7491w7497w7498w7499w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7481w7487w7488w7489w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7471w7477w7478w7479w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7461w7467w7468w7469w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7451w7457w7458w7459w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7441w7447w7448w7449w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7431w7437w7438w7439w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7421w7427w7428w7429w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7411w7417w7418w7419w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7401w7407w7408w7409w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7391w7397w7398w7399w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7381w7387w7388w7389w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7371w7377w7378w7379w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7361w7367w7368w7369w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7351w7357w7358w7359w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7341w7347w7348w7349w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7331w7337w7338w7339w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7321w7327w7328w7329w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7311w7317w7318w7319w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7301w7307w7308w7309w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7291w7297w7298w7299w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7281w7287w7288w7289w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7271w7277w7278w7279w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7261w7267w7268w7269w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7251w7257w7258w7259w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7241w7247w7248w7249w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7231w7237w7238w7239w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7221w7227w7228w7229w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7211w7217w7218w7219w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7201w7207w7208w7209w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7191w7197w7198w7199w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7181w7187w7188w7189w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7171w7177w7178w7179w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7161w7167w7168w7169w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7151w7157w7158w7159w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7141w7147w7148w7149w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7131w7137w7138w7139w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7121w7127w7128w7129w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7111w7117w7118w7119w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7101w7107w7108w7109w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7091w7097w7098w7099w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7081w7087w7088w7089w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7071w7077w7078w7079w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7061w7067w7068w7069w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7051w7057w7058w7059w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7041w7047w7048w7049w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7031w7037w7038w7039w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7021w7027w7028w7029w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7011w7017w7018w7019w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range7001w7007w7008w7009w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6991w6997w6998w6999w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6981w6987w6988w6989w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6971w6977w6978w6979w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6961w6967w6968w6969w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6951w6957w6958w6959w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6941w6947w6948w6949w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6931w6937w6938w6939w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6921w6927w6928w6929w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6911w6917w6918w6919w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6901w6907w6908w6909w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6891w6897w6898w6899w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6881w6887w6888w6889w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6871w6877w6878w6879w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6861w6867w6868w6869w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6851w6857w6858w6859w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6841w6847w6848w6849w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6831w6837w6838w6839w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6821w6827w6828w6829w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6811w6817w6818w6819w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6801w6807w6808w6809w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6791w6797w6798w6799w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6781w6787w6788w6789w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6771w6777w6778w6779w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6761w6767w6768w6769w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6751w6757w6758w6759w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6741w6747w6748w6749w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6731w6737w6738w6739w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6721w6727w6728w6729w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6711w6717w6718w6719w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6701w6707w6708w6709w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6691w6697w6698w6699w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6681w6687w6688w6689w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6671w6677w6678w6679w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6661w6667w6668w6669w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6651w6657w6658w6659w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6641w6647w6648w6649w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6631w6637w6638w6639w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector2_range6619w6626w6627w6628w);
	car_one_adj <= ( car_one(90 DOWNTO 0) & "1");
	car_two <= ( wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8549w8555w8556w8557w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8538w8544w8545w8546w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8527w8533w8534w8535w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8516w8522w8523w8524w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8505w8511w8512w8513w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8494w8500w8501w8502w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8483w8489w8490w8491w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8472w8478w8479w8480w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8461w8467w8468w8469w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8450w8456w8457w8458w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8439w8445w8446w8447w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8428w8434w8435w8436w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8417w8423w8424w8425w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8406w8412w8413w8414w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8395w8401w8402w8403w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8384w8390w8391w8392w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8373w8379w8380w8381w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8362w8368w8369w8370w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8351w8357w8358w8359w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8340w8346w8347w8348w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8329w8335w8336w8337w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8318w8324w8325w8326w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8307w8313w8314w8315w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8296w8302w8303w8304w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8285w8291w8292w8293w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8274w8280w8281w8282w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8263w8269w8270w8271w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8252w8258w8259w8260w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8241w8247w8248w8249w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8230w8236w8237w8238w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8219w8225w8226w8227w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8208w8214w8215w8216w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8197w8203w8204w8205w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8186w8192w8193w8194w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8175w8181w8182w8183w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8164w8170w8171w8172w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8153w8159w8160w8161w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8142w8148w8149w8150w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8131w8137w8138w8139w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8120w8126w8127w8128w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8109w8115w8116w8117w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8098w8104w8105w8106w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8087w8093w8094w8095w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8076w8082w8083w8084w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8065w8071w8072w8073w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8054w8060w8061w8062w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8043w8049w8050w8051w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8032w8038w8039w8040w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8021w8027w8028w8029w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range8010w8016w8017w8018w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7999w8005w8006w8007w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7988w7994w7995w7996w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7977w7983w7984w7985w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7966w7972w7973w7974w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7955w7961w7962w7963w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7944w7950w7951w7952w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7933w7939w7940w7941w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7922w7928w7929w7930w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7911w7917w7918w7919w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7900w7906w7907w7908w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7889w7895w7896w7897w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7878w7884w7885w7886w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7867w7873w7874w7875w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7856w7862w7863w7864w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7845w7851w7852w7853w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7834w7840w7841w7842w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7823w7829w7830w7831w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7812w7818w7819w7820w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7801w7807w7808w7809w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7790w7796w7797w7798w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7779w7785w7786w7787w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7768w7774w7775w7776w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7757w7763w7764w7765w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7746w7752w7753w7754w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7735w7741w7742w7743w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7724w7730w7731w7732w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7713w7719w7720w7721w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7702w7708w7709w7710w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7691w7697w7698w7699w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7680w7686w7687w7688w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7669w7675w7676w7677w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7658w7664w7665w7666w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7647w7653w7654w7655w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7636w7642w7643w7644w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7625w7631w7632w7633w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7614w7620w7621w7622w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7603w7609w7610w7611w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7592w7598w7599w7600w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7581w7587w7588w7589w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7570w7576w7577w7578w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7559w7565w7566w7567w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_lg_w_vector1_range7546w7553w7554w7555w);
	car_two_adj <= ( car_two(90 DOWNTO 0) & "1");
	car_two_wo <= car_two_adj_reg0;
	lowest_bits_wi <= lsb_prod_wo(30 DOWNTO 0);
	lowest_bits_wo <= lowest_bits_wi_reg2;
	lsb_prod_wi <= wire_lsb_prod_result;
	lsb_prod_wo <= lsb_prod_wi_reg0;
	mid_prod_wi <= wire_mid_prod_result;
	mid_prod_wo <= mid_prod_wi_reg0;
	msb_prod_out <= wire_msb_prod_result;
	msb_prod_wi <= msb_prod_out;
	msb_prod_wo <= msb_prod_wi_reg0;
	neg_lsb <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6250w6251w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6256w6257w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6262w6263w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6268w6269w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6274w6275w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6280w6281w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6286w6287w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6292w6293w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6298w6299w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6304w6305w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6310w6311w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6316w6317w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6322w6323w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6328w6329w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6334w6335w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6340w6341w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6346w6347w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6352w6353w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6358w6359w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6364w6365w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6370w6371w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6376w6377w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6382w6383w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6388w6389w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6394w6395w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6400w6401w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6406w6407w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6412w6413w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6418w6419w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6424w6425w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6430w6431w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6436w6437w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6442w6443w
 & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6448w6449w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6454w6455w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6460w6461w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6466w6467w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6472w6473w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6478w6479w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6484w6485w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6490w6491w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6496w6497w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6502w6503w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6508w6509w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6514w6515w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6520w6521w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6526w6527w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6532w6533w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6538w6539w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6544w6545w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6550w6551w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6556w6557w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6562w6563w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6568w6569w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6574w6575w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6580w6581w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6586w6587w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6592w6593w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6598w6599w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6604w6605w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6610w6611w & wire_tbl1_tbl2_prod_w_lg_w_lsb_prod_wo_range6616w6617w);
	neg_msb <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6253w6254w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6259w6260w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6265w6266w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6271w6272w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6277w6278w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6283w6284w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6289w6290w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6295w6296w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6301w6302w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6307w6308w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6313w6314w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6319w6320w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6325w6326w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6331w6332w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6337w6338w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6343w6344w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6349w6350w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6355w6356w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6361w6362w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6367w6368w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6373w6374w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6379w6380w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6385w6386w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6391w6392w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6397w6398w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6403w6404w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6409w6410w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6415w6416w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6421w6422w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6427w6428w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6433w6434w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6439w6440w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6445w6446w
 & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6451w6452w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6457w6458w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6463w6464w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6469w6470w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6475w6476w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6481w6482w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6487w6488w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6493w6494w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6499w6500w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6505w6506w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6511w6512w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6517w6518w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6523w6524w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6529w6530w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6535w6536w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6541w6542w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6547w6548w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6553w6554w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6559w6560w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6565w6566w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6571w6572w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6577w6578w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6583w6584w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6589w6590w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6595w6596w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6601w6602w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6607w6608w & wire_tbl1_tbl2_prod_w_lg_w_msb_prod_wo_range6613w6614w);
	result <= ( wire_sum_result(90 DOWNTO 0) & lowest_bits_wo);
	sum_one <= ( wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7531w7532w7533w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7521w7522w7523w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7511w7512w7513w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7501w7502w7503w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7491w7492w7493w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7481w7482w7483w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7471w7472w7473w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7461w7462w7463w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7451w7452w7453w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7441w7442w7443w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7431w7432w7433w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7421w7422w7423w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7411w7412w7413w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7401w7402w7403w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7391w7392w7393w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7381w7382w7383w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7371w7372w7373w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7361w7362w7363w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7351w7352w7353w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7341w7342w7343w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7331w7332w7333w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7321w7322w7323w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7311w7312w7313w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7301w7302w7303w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7291w7292w7293w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7281w7282w7283w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7271w7272w7273w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7261w7262w7263w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7251w7252w7253w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7241w7242w7243w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7231w7232w7233w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7221w7222w7223w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7211w7212w7213w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7201w7202w7203w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7191w7192w7193w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7181w7182w7183w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7171w7172w7173w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7161w7162w7163w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7151w7152w7153w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7141w7142w7143w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7131w7132w7133w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7121w7122w7123w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7111w7112w7113w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7101w7102w7103w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7091w7092w7093w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7081w7082w7083w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7071w7072w7073w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7061w7062w7063w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7051w7052w7053w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7041w7042w7043w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7031w7032w7033w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7021w7022w7023w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7011w7012w7013w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range7001w7002w7003w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6991w6992w6993w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6981w6982w6983w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6971w6972w6973w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6961w6962w6963w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6951w6952w6953w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6941w6942w6943w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6931w6932w6933w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6921w6922w6923w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6911w6912w6913w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6901w6902w6903w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6891w6892w6893w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6881w6882w6883w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6871w6872w6873w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6861w6862w6863w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6851w6852w6853w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6841w6842w6843w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6831w6832w6833w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6821w6822w6823w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6811w6812w6813w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6801w6802w6803w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6791w6792w6793w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6781w6782w6783w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6771w6772w6773w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6761w6762w6763w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6751w6752w6753w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6741w6742w6743w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6731w6732w6733w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6721w6722w6723w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6711w6712w6713w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6701w6702w6703w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6691w6692w6693w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6681w6682w6683w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6671w6672w6673w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6661w6662w6663w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6651w6652w6653w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6641w6642w6643w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6631w6632w6633w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector2_range6619w6620w6621w);
	sum_two <= ( wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8549w8550w8551w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8538w8539w8540w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8527w8528w8529w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8516w8517w8518w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8505w8506w8507w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8494w8495w8496w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8483w8484w8485w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8472w8473w8474w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8461w8462w8463w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8450w8451w8452w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8439w8440w8441w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8428w8429w8430w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8417w8418w8419w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8406w8407w8408w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8395w8396w8397w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8384w8385w8386w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8373w8374w8375w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8362w8363w8364w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8351w8352w8353w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8340w8341w8342w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8329w8330w8331w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8318w8319w8320w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8307w8308w8309w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8296w8297w8298w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8285w8286w8287w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8274w8275w8276w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8263w8264w8265w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8252w8253w8254w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8241w8242w8243w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8230w8231w8232w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8219w8220w8221w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8208w8209w8210w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8197w8198w8199w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8186w8187w8188w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8175w8176w8177w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8164w8165w8166w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8153w8154w8155w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8142w8143w8144w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8131w8132w8133w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8120w8121w8122w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8109w8110w8111w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8098w8099w8100w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8087w8088w8089w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8076w8077w8078w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8065w8066w8067w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8054w8055w8056w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8043w8044w8045w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8032w8033w8034w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8021w8022w8023w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range8010w8011w8012w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7999w8000w8001w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7988w7989w7990w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7977w7978w7979w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7966w7967w7968w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7955w7956w7957w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7944w7945w7946w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7933w7934w7935w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7922w7923w7924w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7911w7912w7913w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7900w7901w7902w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7889w7890w7891w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7878w7879w7880w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7867w7868w7869w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7856w7857w7858w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7845w7846w7847w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7834w7835w7836w
 & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7823w7824w7825w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7812w7813w7814w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7801w7802w7803w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7790w7791w7792w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7779w7780w7781w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7768w7769w7770w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7757w7758w7759w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7746w7747w7748w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7735w7736w7737w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7724w7725w7726w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7713w7714w7715w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7702w7703w7704w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7691w7692w7693w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7680w7681w7682w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7669w7670w7671w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7658w7659w7660w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7647w7648w7649w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7636w7637w7638w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7625w7626w7627w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7614w7615w7616w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7603w7604w7605w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7592w7593w7594w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7581w7582w7583w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7570w7571w7572w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7559w7560w7561w & wire_tbl1_tbl2_prod_w_lg_w_lg_w_vector1_range7546w7547w7548w);
	sum_two_wo <= sum_two_reg0;
	vector1 <= ( msb_prod_wo & lsb_prod_wo(61 DOWNTO 31));
	vector2 <= ( "0000000000000000000000000000" & mid_prod_wo);
	wire_a <= dataa;
	wire_b <= datab;
	wire_tbl1_tbl2_prod_w_car_one_adj_range7544w(0) <= car_one_adj(0);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7657w(0) <= car_one_adj(10);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7668w(0) <= car_one_adj(11);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7679w(0) <= car_one_adj(12);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7690w(0) <= car_one_adj(13);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7701w(0) <= car_one_adj(14);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7712w(0) <= car_one_adj(15);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7723w(0) <= car_one_adj(16);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7734w(0) <= car_one_adj(17);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7745w(0) <= car_one_adj(18);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7756w(0) <= car_one_adj(19);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7558w(0) <= car_one_adj(1);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7767w(0) <= car_one_adj(20);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7778w(0) <= car_one_adj(21);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7789w(0) <= car_one_adj(22);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7800w(0) <= car_one_adj(23);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7811w(0) <= car_one_adj(24);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7822w(0) <= car_one_adj(25);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7833w(0) <= car_one_adj(26);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7844w(0) <= car_one_adj(27);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7855w(0) <= car_one_adj(28);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7866w(0) <= car_one_adj(29);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7569w(0) <= car_one_adj(2);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7877w(0) <= car_one_adj(30);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7888w(0) <= car_one_adj(31);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7899w(0) <= car_one_adj(32);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7910w(0) <= car_one_adj(33);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7921w(0) <= car_one_adj(34);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7932w(0) <= car_one_adj(35);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7943w(0) <= car_one_adj(36);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7954w(0) <= car_one_adj(37);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7965w(0) <= car_one_adj(38);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7976w(0) <= car_one_adj(39);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7580w(0) <= car_one_adj(3);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7987w(0) <= car_one_adj(40);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7998w(0) <= car_one_adj(41);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8009w(0) <= car_one_adj(42);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8020w(0) <= car_one_adj(43);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8031w(0) <= car_one_adj(44);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8042w(0) <= car_one_adj(45);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8053w(0) <= car_one_adj(46);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8064w(0) <= car_one_adj(47);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8075w(0) <= car_one_adj(48);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8086w(0) <= car_one_adj(49);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7591w(0) <= car_one_adj(4);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8097w(0) <= car_one_adj(50);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8108w(0) <= car_one_adj(51);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8119w(0) <= car_one_adj(52);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8130w(0) <= car_one_adj(53);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8141w(0) <= car_one_adj(54);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8152w(0) <= car_one_adj(55);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8163w(0) <= car_one_adj(56);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8174w(0) <= car_one_adj(57);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8185w(0) <= car_one_adj(58);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8196w(0) <= car_one_adj(59);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7602w(0) <= car_one_adj(5);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8207w(0) <= car_one_adj(60);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8218w(0) <= car_one_adj(61);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8229w(0) <= car_one_adj(62);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8240w(0) <= car_one_adj(63);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8251w(0) <= car_one_adj(64);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8262w(0) <= car_one_adj(65);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8273w(0) <= car_one_adj(66);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8284w(0) <= car_one_adj(67);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8295w(0) <= car_one_adj(68);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8306w(0) <= car_one_adj(69);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7613w(0) <= car_one_adj(6);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8317w(0) <= car_one_adj(70);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8328w(0) <= car_one_adj(71);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8339w(0) <= car_one_adj(72);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8350w(0) <= car_one_adj(73);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8361w(0) <= car_one_adj(74);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8372w(0) <= car_one_adj(75);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8383w(0) <= car_one_adj(76);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8394w(0) <= car_one_adj(77);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8405w(0) <= car_one_adj(78);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8416w(0) <= car_one_adj(79);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7624w(0) <= car_one_adj(7);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8427w(0) <= car_one_adj(80);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8438w(0) <= car_one_adj(81);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8449w(0) <= car_one_adj(82);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8460w(0) <= car_one_adj(83);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8471w(0) <= car_one_adj(84);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8482w(0) <= car_one_adj(85);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8493w(0) <= car_one_adj(86);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8504w(0) <= car_one_adj(87);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8515w(0) <= car_one_adj(88);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8526w(0) <= car_one_adj(89);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7635w(0) <= car_one_adj(8);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8537w(0) <= car_one_adj(90);
	wire_tbl1_tbl2_prod_w_car_one_adj_range8548w(0) <= car_one_adj(91);
	wire_tbl1_tbl2_prod_w_car_one_adj_range7646w(0) <= car_one_adj(9);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6616w(0) <= lsb_prod_wo(0);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6556w(0) <= lsb_prod_wo(10);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6550w(0) <= lsb_prod_wo(11);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6544w(0) <= lsb_prod_wo(12);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6538w(0) <= lsb_prod_wo(13);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6532w(0) <= lsb_prod_wo(14);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6526w(0) <= lsb_prod_wo(15);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6520w(0) <= lsb_prod_wo(16);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6514w(0) <= lsb_prod_wo(17);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6508w(0) <= lsb_prod_wo(18);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6502w(0) <= lsb_prod_wo(19);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6610w(0) <= lsb_prod_wo(1);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6496w(0) <= lsb_prod_wo(20);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6490w(0) <= lsb_prod_wo(21);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6484w(0) <= lsb_prod_wo(22);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6478w(0) <= lsb_prod_wo(23);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6472w(0) <= lsb_prod_wo(24);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6466w(0) <= lsb_prod_wo(25);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6460w(0) <= lsb_prod_wo(26);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6454w(0) <= lsb_prod_wo(27);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6448w(0) <= lsb_prod_wo(28);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6442w(0) <= lsb_prod_wo(29);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6604w(0) <= lsb_prod_wo(2);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6436w(0) <= lsb_prod_wo(30);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6430w(0) <= lsb_prod_wo(31);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6424w(0) <= lsb_prod_wo(32);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6418w(0) <= lsb_prod_wo(33);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6412w(0) <= lsb_prod_wo(34);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6406w(0) <= lsb_prod_wo(35);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6400w(0) <= lsb_prod_wo(36);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6394w(0) <= lsb_prod_wo(37);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6388w(0) <= lsb_prod_wo(38);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6382w(0) <= lsb_prod_wo(39);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6598w(0) <= lsb_prod_wo(3);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6376w(0) <= lsb_prod_wo(40);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6370w(0) <= lsb_prod_wo(41);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6364w(0) <= lsb_prod_wo(42);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6358w(0) <= lsb_prod_wo(43);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6352w(0) <= lsb_prod_wo(44);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6346w(0) <= lsb_prod_wo(45);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6340w(0) <= lsb_prod_wo(46);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6334w(0) <= lsb_prod_wo(47);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6328w(0) <= lsb_prod_wo(48);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6322w(0) <= lsb_prod_wo(49);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6592w(0) <= lsb_prod_wo(4);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6316w(0) <= lsb_prod_wo(50);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6310w(0) <= lsb_prod_wo(51);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6304w(0) <= lsb_prod_wo(52);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6298w(0) <= lsb_prod_wo(53);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6292w(0) <= lsb_prod_wo(54);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6286w(0) <= lsb_prod_wo(55);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6280w(0) <= lsb_prod_wo(56);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6274w(0) <= lsb_prod_wo(57);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6268w(0) <= lsb_prod_wo(58);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6262w(0) <= lsb_prod_wo(59);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6586w(0) <= lsb_prod_wo(5);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6256w(0) <= lsb_prod_wo(60);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6250w(0) <= lsb_prod_wo(61);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6580w(0) <= lsb_prod_wo(6);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6574w(0) <= lsb_prod_wo(7);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6568w(0) <= lsb_prod_wo(8);
	wire_tbl1_tbl2_prod_w_lsb_prod_wo_range6562w(0) <= lsb_prod_wo(9);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6613w(0) <= msb_prod_wo(0);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6553w(0) <= msb_prod_wo(10);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6547w(0) <= msb_prod_wo(11);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6541w(0) <= msb_prod_wo(12);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6535w(0) <= msb_prod_wo(13);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6529w(0) <= msb_prod_wo(14);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6523w(0) <= msb_prod_wo(15);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6517w(0) <= msb_prod_wo(16);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6511w(0) <= msb_prod_wo(17);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6505w(0) <= msb_prod_wo(18);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6499w(0) <= msb_prod_wo(19);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6607w(0) <= msb_prod_wo(1);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6493w(0) <= msb_prod_wo(20);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6487w(0) <= msb_prod_wo(21);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6481w(0) <= msb_prod_wo(22);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6475w(0) <= msb_prod_wo(23);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6469w(0) <= msb_prod_wo(24);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6463w(0) <= msb_prod_wo(25);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6457w(0) <= msb_prod_wo(26);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6451w(0) <= msb_prod_wo(27);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6445w(0) <= msb_prod_wo(28);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6439w(0) <= msb_prod_wo(29);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6601w(0) <= msb_prod_wo(2);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6433w(0) <= msb_prod_wo(30);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6427w(0) <= msb_prod_wo(31);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6421w(0) <= msb_prod_wo(32);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6415w(0) <= msb_prod_wo(33);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6409w(0) <= msb_prod_wo(34);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6403w(0) <= msb_prod_wo(35);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6397w(0) <= msb_prod_wo(36);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6391w(0) <= msb_prod_wo(37);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6385w(0) <= msb_prod_wo(38);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6379w(0) <= msb_prod_wo(39);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6595w(0) <= msb_prod_wo(3);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6373w(0) <= msb_prod_wo(40);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6367w(0) <= msb_prod_wo(41);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6361w(0) <= msb_prod_wo(42);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6355w(0) <= msb_prod_wo(43);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6349w(0) <= msb_prod_wo(44);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6343w(0) <= msb_prod_wo(45);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6337w(0) <= msb_prod_wo(46);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6331w(0) <= msb_prod_wo(47);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6325w(0) <= msb_prod_wo(48);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6319w(0) <= msb_prod_wo(49);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6589w(0) <= msb_prod_wo(4);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6313w(0) <= msb_prod_wo(50);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6307w(0) <= msb_prod_wo(51);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6301w(0) <= msb_prod_wo(52);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6295w(0) <= msb_prod_wo(53);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6289w(0) <= msb_prod_wo(54);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6283w(0) <= msb_prod_wo(55);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6277w(0) <= msb_prod_wo(56);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6271w(0) <= msb_prod_wo(57);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6265w(0) <= msb_prod_wo(58);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6259w(0) <= msb_prod_wo(59);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6583w(0) <= msb_prod_wo(5);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6253w(0) <= msb_prod_wo(60);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6577w(0) <= msb_prod_wo(6);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6571w(0) <= msb_prod_wo(7);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6565w(0) <= msb_prod_wo(8);
	wire_tbl1_tbl2_prod_w_msb_prod_wo_range6559w(0) <= msb_prod_wo(9);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6618w(0) <= neg_lsb(0);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6558w(0) <= neg_lsb(10);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6552w(0) <= neg_lsb(11);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6546w(0) <= neg_lsb(12);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6540w(0) <= neg_lsb(13);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6534w(0) <= neg_lsb(14);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6528w(0) <= neg_lsb(15);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6522w(0) <= neg_lsb(16);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6516w(0) <= neg_lsb(17);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6510w(0) <= neg_lsb(18);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6504w(0) <= neg_lsb(19);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6612w(0) <= neg_lsb(1);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6498w(0) <= neg_lsb(20);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6492w(0) <= neg_lsb(21);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6486w(0) <= neg_lsb(22);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6480w(0) <= neg_lsb(23);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6474w(0) <= neg_lsb(24);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6468w(0) <= neg_lsb(25);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6462w(0) <= neg_lsb(26);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6456w(0) <= neg_lsb(27);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6450w(0) <= neg_lsb(28);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6444w(0) <= neg_lsb(29);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6606w(0) <= neg_lsb(2);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6438w(0) <= neg_lsb(30);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6432w(0) <= neg_lsb(31);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6426w(0) <= neg_lsb(32);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6420w(0) <= neg_lsb(33);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6414w(0) <= neg_lsb(34);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6408w(0) <= neg_lsb(35);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6402w(0) <= neg_lsb(36);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6396w(0) <= neg_lsb(37);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6390w(0) <= neg_lsb(38);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6384w(0) <= neg_lsb(39);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6600w(0) <= neg_lsb(3);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6378w(0) <= neg_lsb(40);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6372w(0) <= neg_lsb(41);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6366w(0) <= neg_lsb(42);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6360w(0) <= neg_lsb(43);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6354w(0) <= neg_lsb(44);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6348w(0) <= neg_lsb(45);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6342w(0) <= neg_lsb(46);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6336w(0) <= neg_lsb(47);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6330w(0) <= neg_lsb(48);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6324w(0) <= neg_lsb(49);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6594w(0) <= neg_lsb(4);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6318w(0) <= neg_lsb(50);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6312w(0) <= neg_lsb(51);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6306w(0) <= neg_lsb(52);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6300w(0) <= neg_lsb(53);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6294w(0) <= neg_lsb(54);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6288w(0) <= neg_lsb(55);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6282w(0) <= neg_lsb(56);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6276w(0) <= neg_lsb(57);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6270w(0) <= neg_lsb(58);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6264w(0) <= neg_lsb(59);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6588w(0) <= neg_lsb(5);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6258w(0) <= neg_lsb(60);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6252w(0) <= neg_lsb(61);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6246w(0) <= neg_lsb(62);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6242w(0) <= neg_lsb(63);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6238w(0) <= neg_lsb(64);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6234w(0) <= neg_lsb(65);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6230w(0) <= neg_lsb(66);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6226w(0) <= neg_lsb(67);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6222w(0) <= neg_lsb(68);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6218w(0) <= neg_lsb(69);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6582w(0) <= neg_lsb(6);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6214w(0) <= neg_lsb(70);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6210w(0) <= neg_lsb(71);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6206w(0) <= neg_lsb(72);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6202w(0) <= neg_lsb(73);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6198w(0) <= neg_lsb(74);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6194w(0) <= neg_lsb(75);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6190w(0) <= neg_lsb(76);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6186w(0) <= neg_lsb(77);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6182w(0) <= neg_lsb(78);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6178w(0) <= neg_lsb(79);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6576w(0) <= neg_lsb(7);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6174w(0) <= neg_lsb(80);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6170w(0) <= neg_lsb(81);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6166w(0) <= neg_lsb(82);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6162w(0) <= neg_lsb(83);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6158w(0) <= neg_lsb(84);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6154w(0) <= neg_lsb(85);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6150w(0) <= neg_lsb(86);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6146w(0) <= neg_lsb(87);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6142w(0) <= neg_lsb(88);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6138w(0) <= neg_lsb(89);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6570w(0) <= neg_lsb(8);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6134w(0) <= neg_lsb(90);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6129w(0) <= neg_lsb(91);
	wire_tbl1_tbl2_prod_w_neg_lsb_range6564w(0) <= neg_lsb(9);
	wire_tbl1_tbl2_prod_w_neg_msb_range6615w(0) <= neg_msb(0);
	wire_tbl1_tbl2_prod_w_neg_msb_range6555w(0) <= neg_msb(10);
	wire_tbl1_tbl2_prod_w_neg_msb_range6549w(0) <= neg_msb(11);
	wire_tbl1_tbl2_prod_w_neg_msb_range6543w(0) <= neg_msb(12);
	wire_tbl1_tbl2_prod_w_neg_msb_range6537w(0) <= neg_msb(13);
	wire_tbl1_tbl2_prod_w_neg_msb_range6531w(0) <= neg_msb(14);
	wire_tbl1_tbl2_prod_w_neg_msb_range6525w(0) <= neg_msb(15);
	wire_tbl1_tbl2_prod_w_neg_msb_range6519w(0) <= neg_msb(16);
	wire_tbl1_tbl2_prod_w_neg_msb_range6513w(0) <= neg_msb(17);
	wire_tbl1_tbl2_prod_w_neg_msb_range6507w(0) <= neg_msb(18);
	wire_tbl1_tbl2_prod_w_neg_msb_range6501w(0) <= neg_msb(19);
	wire_tbl1_tbl2_prod_w_neg_msb_range6609w(0) <= neg_msb(1);
	wire_tbl1_tbl2_prod_w_neg_msb_range6495w(0) <= neg_msb(20);
	wire_tbl1_tbl2_prod_w_neg_msb_range6489w(0) <= neg_msb(21);
	wire_tbl1_tbl2_prod_w_neg_msb_range6483w(0) <= neg_msb(22);
	wire_tbl1_tbl2_prod_w_neg_msb_range6477w(0) <= neg_msb(23);
	wire_tbl1_tbl2_prod_w_neg_msb_range6471w(0) <= neg_msb(24);
	wire_tbl1_tbl2_prod_w_neg_msb_range6465w(0) <= neg_msb(25);
	wire_tbl1_tbl2_prod_w_neg_msb_range6459w(0) <= neg_msb(26);
	wire_tbl1_tbl2_prod_w_neg_msb_range6453w(0) <= neg_msb(27);
	wire_tbl1_tbl2_prod_w_neg_msb_range6447w(0) <= neg_msb(28);
	wire_tbl1_tbl2_prod_w_neg_msb_range6441w(0) <= neg_msb(29);
	wire_tbl1_tbl2_prod_w_neg_msb_range6603w(0) <= neg_msb(2);
	wire_tbl1_tbl2_prod_w_neg_msb_range6435w(0) <= neg_msb(30);
	wire_tbl1_tbl2_prod_w_neg_msb_range6429w(0) <= neg_msb(31);
	wire_tbl1_tbl2_prod_w_neg_msb_range6423w(0) <= neg_msb(32);
	wire_tbl1_tbl2_prod_w_neg_msb_range6417w(0) <= neg_msb(33);
	wire_tbl1_tbl2_prod_w_neg_msb_range6411w(0) <= neg_msb(34);
	wire_tbl1_tbl2_prod_w_neg_msb_range6405w(0) <= neg_msb(35);
	wire_tbl1_tbl2_prod_w_neg_msb_range6399w(0) <= neg_msb(36);
	wire_tbl1_tbl2_prod_w_neg_msb_range6393w(0) <= neg_msb(37);
	wire_tbl1_tbl2_prod_w_neg_msb_range6387w(0) <= neg_msb(38);
	wire_tbl1_tbl2_prod_w_neg_msb_range6381w(0) <= neg_msb(39);
	wire_tbl1_tbl2_prod_w_neg_msb_range6597w(0) <= neg_msb(3);
	wire_tbl1_tbl2_prod_w_neg_msb_range6375w(0) <= neg_msb(40);
	wire_tbl1_tbl2_prod_w_neg_msb_range6369w(0) <= neg_msb(41);
	wire_tbl1_tbl2_prod_w_neg_msb_range6363w(0) <= neg_msb(42);
	wire_tbl1_tbl2_prod_w_neg_msb_range6357w(0) <= neg_msb(43);
	wire_tbl1_tbl2_prod_w_neg_msb_range6351w(0) <= neg_msb(44);
	wire_tbl1_tbl2_prod_w_neg_msb_range6345w(0) <= neg_msb(45);
	wire_tbl1_tbl2_prod_w_neg_msb_range6339w(0) <= neg_msb(46);
	wire_tbl1_tbl2_prod_w_neg_msb_range6333w(0) <= neg_msb(47);
	wire_tbl1_tbl2_prod_w_neg_msb_range6327w(0) <= neg_msb(48);
	wire_tbl1_tbl2_prod_w_neg_msb_range6321w(0) <= neg_msb(49);
	wire_tbl1_tbl2_prod_w_neg_msb_range6591w(0) <= neg_msb(4);
	wire_tbl1_tbl2_prod_w_neg_msb_range6315w(0) <= neg_msb(50);
	wire_tbl1_tbl2_prod_w_neg_msb_range6309w(0) <= neg_msb(51);
	wire_tbl1_tbl2_prod_w_neg_msb_range6303w(0) <= neg_msb(52);
	wire_tbl1_tbl2_prod_w_neg_msb_range6297w(0) <= neg_msb(53);
	wire_tbl1_tbl2_prod_w_neg_msb_range6291w(0) <= neg_msb(54);
	wire_tbl1_tbl2_prod_w_neg_msb_range6285w(0) <= neg_msb(55);
	wire_tbl1_tbl2_prod_w_neg_msb_range6279w(0) <= neg_msb(56);
	wire_tbl1_tbl2_prod_w_neg_msb_range6273w(0) <= neg_msb(57);
	wire_tbl1_tbl2_prod_w_neg_msb_range6267w(0) <= neg_msb(58);
	wire_tbl1_tbl2_prod_w_neg_msb_range6261w(0) <= neg_msb(59);
	wire_tbl1_tbl2_prod_w_neg_msb_range6585w(0) <= neg_msb(5);
	wire_tbl1_tbl2_prod_w_neg_msb_range6255w(0) <= neg_msb(60);
	wire_tbl1_tbl2_prod_w_neg_msb_range6248w(0) <= neg_msb(61);
	wire_tbl1_tbl2_prod_w_neg_msb_range6244w(0) <= neg_msb(62);
	wire_tbl1_tbl2_prod_w_neg_msb_range6240w(0) <= neg_msb(63);
	wire_tbl1_tbl2_prod_w_neg_msb_range6236w(0) <= neg_msb(64);
	wire_tbl1_tbl2_prod_w_neg_msb_range6232w(0) <= neg_msb(65);
	wire_tbl1_tbl2_prod_w_neg_msb_range6228w(0) <= neg_msb(66);
	wire_tbl1_tbl2_prod_w_neg_msb_range6224w(0) <= neg_msb(67);
	wire_tbl1_tbl2_prod_w_neg_msb_range6220w(0) <= neg_msb(68);
	wire_tbl1_tbl2_prod_w_neg_msb_range6216w(0) <= neg_msb(69);
	wire_tbl1_tbl2_prod_w_neg_msb_range6579w(0) <= neg_msb(6);
	wire_tbl1_tbl2_prod_w_neg_msb_range6212w(0) <= neg_msb(70);
	wire_tbl1_tbl2_prod_w_neg_msb_range6208w(0) <= neg_msb(71);
	wire_tbl1_tbl2_prod_w_neg_msb_range6204w(0) <= neg_msb(72);
	wire_tbl1_tbl2_prod_w_neg_msb_range6200w(0) <= neg_msb(73);
	wire_tbl1_tbl2_prod_w_neg_msb_range6196w(0) <= neg_msb(74);
	wire_tbl1_tbl2_prod_w_neg_msb_range6192w(0) <= neg_msb(75);
	wire_tbl1_tbl2_prod_w_neg_msb_range6188w(0) <= neg_msb(76);
	wire_tbl1_tbl2_prod_w_neg_msb_range6184w(0) <= neg_msb(77);
	wire_tbl1_tbl2_prod_w_neg_msb_range6180w(0) <= neg_msb(78);
	wire_tbl1_tbl2_prod_w_neg_msb_range6176w(0) <= neg_msb(79);
	wire_tbl1_tbl2_prod_w_neg_msb_range6573w(0) <= neg_msb(7);
	wire_tbl1_tbl2_prod_w_neg_msb_range6172w(0) <= neg_msb(80);
	wire_tbl1_tbl2_prod_w_neg_msb_range6168w(0) <= neg_msb(81);
	wire_tbl1_tbl2_prod_w_neg_msb_range6164w(0) <= neg_msb(82);
	wire_tbl1_tbl2_prod_w_neg_msb_range6160w(0) <= neg_msb(83);
	wire_tbl1_tbl2_prod_w_neg_msb_range6156w(0) <= neg_msb(84);
	wire_tbl1_tbl2_prod_w_neg_msb_range6152w(0) <= neg_msb(85);
	wire_tbl1_tbl2_prod_w_neg_msb_range6148w(0) <= neg_msb(86);
	wire_tbl1_tbl2_prod_w_neg_msb_range6144w(0) <= neg_msb(87);
	wire_tbl1_tbl2_prod_w_neg_msb_range6140w(0) <= neg_msb(88);
	wire_tbl1_tbl2_prod_w_neg_msb_range6136w(0) <= neg_msb(89);
	wire_tbl1_tbl2_prod_w_neg_msb_range6567w(0) <= neg_msb(8);
	wire_tbl1_tbl2_prod_w_neg_msb_range6132w(0) <= neg_msb(90);
	wire_tbl1_tbl2_prod_w_neg_msb_range6126w(0) <= neg_msb(91);
	wire_tbl1_tbl2_prod_w_neg_msb_range6561w(0) <= neg_msb(9);
	wire_tbl1_tbl2_prod_w_sum_one_range6622w(0) <= sum_one(0);
	wire_tbl1_tbl2_prod_w_sum_one_range6724w(0) <= sum_one(10);
	wire_tbl1_tbl2_prod_w_sum_one_range6734w(0) <= sum_one(11);
	wire_tbl1_tbl2_prod_w_sum_one_range6744w(0) <= sum_one(12);
	wire_tbl1_tbl2_prod_w_sum_one_range6754w(0) <= sum_one(13);
	wire_tbl1_tbl2_prod_w_sum_one_range6764w(0) <= sum_one(14);
	wire_tbl1_tbl2_prod_w_sum_one_range6774w(0) <= sum_one(15);
	wire_tbl1_tbl2_prod_w_sum_one_range6784w(0) <= sum_one(16);
	wire_tbl1_tbl2_prod_w_sum_one_range6794w(0) <= sum_one(17);
	wire_tbl1_tbl2_prod_w_sum_one_range6804w(0) <= sum_one(18);
	wire_tbl1_tbl2_prod_w_sum_one_range6814w(0) <= sum_one(19);
	wire_tbl1_tbl2_prod_w_sum_one_range6634w(0) <= sum_one(1);
	wire_tbl1_tbl2_prod_w_sum_one_range6824w(0) <= sum_one(20);
	wire_tbl1_tbl2_prod_w_sum_one_range6834w(0) <= sum_one(21);
	wire_tbl1_tbl2_prod_w_sum_one_range6844w(0) <= sum_one(22);
	wire_tbl1_tbl2_prod_w_sum_one_range6854w(0) <= sum_one(23);
	wire_tbl1_tbl2_prod_w_sum_one_range6864w(0) <= sum_one(24);
	wire_tbl1_tbl2_prod_w_sum_one_range6874w(0) <= sum_one(25);
	wire_tbl1_tbl2_prod_w_sum_one_range6884w(0) <= sum_one(26);
	wire_tbl1_tbl2_prod_w_sum_one_range6894w(0) <= sum_one(27);
	wire_tbl1_tbl2_prod_w_sum_one_range6904w(0) <= sum_one(28);
	wire_tbl1_tbl2_prod_w_sum_one_range6914w(0) <= sum_one(29);
	wire_tbl1_tbl2_prod_w_sum_one_range6644w(0) <= sum_one(2);
	wire_tbl1_tbl2_prod_w_sum_one_range6924w(0) <= sum_one(30);
	wire_tbl1_tbl2_prod_w_sum_one_range6934w(0) <= sum_one(31);
	wire_tbl1_tbl2_prod_w_sum_one_range6944w(0) <= sum_one(32);
	wire_tbl1_tbl2_prod_w_sum_one_range6954w(0) <= sum_one(33);
	wire_tbl1_tbl2_prod_w_sum_one_range6964w(0) <= sum_one(34);
	wire_tbl1_tbl2_prod_w_sum_one_range6974w(0) <= sum_one(35);
	wire_tbl1_tbl2_prod_w_sum_one_range6984w(0) <= sum_one(36);
	wire_tbl1_tbl2_prod_w_sum_one_range6994w(0) <= sum_one(37);
	wire_tbl1_tbl2_prod_w_sum_one_range7004w(0) <= sum_one(38);
	wire_tbl1_tbl2_prod_w_sum_one_range7014w(0) <= sum_one(39);
	wire_tbl1_tbl2_prod_w_sum_one_range6654w(0) <= sum_one(3);
	wire_tbl1_tbl2_prod_w_sum_one_range7024w(0) <= sum_one(40);
	wire_tbl1_tbl2_prod_w_sum_one_range7034w(0) <= sum_one(41);
	wire_tbl1_tbl2_prod_w_sum_one_range7044w(0) <= sum_one(42);
	wire_tbl1_tbl2_prod_w_sum_one_range7054w(0) <= sum_one(43);
	wire_tbl1_tbl2_prod_w_sum_one_range7064w(0) <= sum_one(44);
	wire_tbl1_tbl2_prod_w_sum_one_range7074w(0) <= sum_one(45);
	wire_tbl1_tbl2_prod_w_sum_one_range7084w(0) <= sum_one(46);
	wire_tbl1_tbl2_prod_w_sum_one_range7094w(0) <= sum_one(47);
	wire_tbl1_tbl2_prod_w_sum_one_range7104w(0) <= sum_one(48);
	wire_tbl1_tbl2_prod_w_sum_one_range7114w(0) <= sum_one(49);
	wire_tbl1_tbl2_prod_w_sum_one_range6664w(0) <= sum_one(4);
	wire_tbl1_tbl2_prod_w_sum_one_range7124w(0) <= sum_one(50);
	wire_tbl1_tbl2_prod_w_sum_one_range7134w(0) <= sum_one(51);
	wire_tbl1_tbl2_prod_w_sum_one_range7144w(0) <= sum_one(52);
	wire_tbl1_tbl2_prod_w_sum_one_range7154w(0) <= sum_one(53);
	wire_tbl1_tbl2_prod_w_sum_one_range7164w(0) <= sum_one(54);
	wire_tbl1_tbl2_prod_w_sum_one_range7174w(0) <= sum_one(55);
	wire_tbl1_tbl2_prod_w_sum_one_range7184w(0) <= sum_one(56);
	wire_tbl1_tbl2_prod_w_sum_one_range7194w(0) <= sum_one(57);
	wire_tbl1_tbl2_prod_w_sum_one_range7204w(0) <= sum_one(58);
	wire_tbl1_tbl2_prod_w_sum_one_range7214w(0) <= sum_one(59);
	wire_tbl1_tbl2_prod_w_sum_one_range6674w(0) <= sum_one(5);
	wire_tbl1_tbl2_prod_w_sum_one_range7224w(0) <= sum_one(60);
	wire_tbl1_tbl2_prod_w_sum_one_range7234w(0) <= sum_one(61);
	wire_tbl1_tbl2_prod_w_sum_one_range7244w(0) <= sum_one(62);
	wire_tbl1_tbl2_prod_w_sum_one_range7254w(0) <= sum_one(63);
	wire_tbl1_tbl2_prod_w_sum_one_range7264w(0) <= sum_one(64);
	wire_tbl1_tbl2_prod_w_sum_one_range7274w(0) <= sum_one(65);
	wire_tbl1_tbl2_prod_w_sum_one_range7284w(0) <= sum_one(66);
	wire_tbl1_tbl2_prod_w_sum_one_range7294w(0) <= sum_one(67);
	wire_tbl1_tbl2_prod_w_sum_one_range7304w(0) <= sum_one(68);
	wire_tbl1_tbl2_prod_w_sum_one_range7314w(0) <= sum_one(69);
	wire_tbl1_tbl2_prod_w_sum_one_range6684w(0) <= sum_one(6);
	wire_tbl1_tbl2_prod_w_sum_one_range7324w(0) <= sum_one(70);
	wire_tbl1_tbl2_prod_w_sum_one_range7334w(0) <= sum_one(71);
	wire_tbl1_tbl2_prod_w_sum_one_range7344w(0) <= sum_one(72);
	wire_tbl1_tbl2_prod_w_sum_one_range7354w(0) <= sum_one(73);
	wire_tbl1_tbl2_prod_w_sum_one_range7364w(0) <= sum_one(74);
	wire_tbl1_tbl2_prod_w_sum_one_range7374w(0) <= sum_one(75);
	wire_tbl1_tbl2_prod_w_sum_one_range7384w(0) <= sum_one(76);
	wire_tbl1_tbl2_prod_w_sum_one_range7394w(0) <= sum_one(77);
	wire_tbl1_tbl2_prod_w_sum_one_range7404w(0) <= sum_one(78);
	wire_tbl1_tbl2_prod_w_sum_one_range7414w(0) <= sum_one(79);
	wire_tbl1_tbl2_prod_w_sum_one_range6694w(0) <= sum_one(7);
	wire_tbl1_tbl2_prod_w_sum_one_range7424w(0) <= sum_one(80);
	wire_tbl1_tbl2_prod_w_sum_one_range7434w(0) <= sum_one(81);
	wire_tbl1_tbl2_prod_w_sum_one_range7444w(0) <= sum_one(82);
	wire_tbl1_tbl2_prod_w_sum_one_range7454w(0) <= sum_one(83);
	wire_tbl1_tbl2_prod_w_sum_one_range7464w(0) <= sum_one(84);
	wire_tbl1_tbl2_prod_w_sum_one_range7474w(0) <= sum_one(85);
	wire_tbl1_tbl2_prod_w_sum_one_range7484w(0) <= sum_one(86);
	wire_tbl1_tbl2_prod_w_sum_one_range7494w(0) <= sum_one(87);
	wire_tbl1_tbl2_prod_w_sum_one_range7504w(0) <= sum_one(88);
	wire_tbl1_tbl2_prod_w_sum_one_range7514w(0) <= sum_one(89);
	wire_tbl1_tbl2_prod_w_sum_one_range6704w(0) <= sum_one(8);
	wire_tbl1_tbl2_prod_w_sum_one_range7524w(0) <= sum_one(90);
	wire_tbl1_tbl2_prod_w_sum_one_range7534w(0) <= sum_one(91);
	wire_tbl1_tbl2_prod_w_sum_one_range6714w(0) <= sum_one(9);
	wire_tbl1_tbl2_prod_w_vector1_range7546w(0) <= vector1(0);
	wire_tbl1_tbl2_prod_w_vector1_range7658w(0) <= vector1(10);
	wire_tbl1_tbl2_prod_w_vector1_range7669w(0) <= vector1(11);
	wire_tbl1_tbl2_prod_w_vector1_range7680w(0) <= vector1(12);
	wire_tbl1_tbl2_prod_w_vector1_range7691w(0) <= vector1(13);
	wire_tbl1_tbl2_prod_w_vector1_range7702w(0) <= vector1(14);
	wire_tbl1_tbl2_prod_w_vector1_range7713w(0) <= vector1(15);
	wire_tbl1_tbl2_prod_w_vector1_range7724w(0) <= vector1(16);
	wire_tbl1_tbl2_prod_w_vector1_range7735w(0) <= vector1(17);
	wire_tbl1_tbl2_prod_w_vector1_range7746w(0) <= vector1(18);
	wire_tbl1_tbl2_prod_w_vector1_range7757w(0) <= vector1(19);
	wire_tbl1_tbl2_prod_w_vector1_range7559w(0) <= vector1(1);
	wire_tbl1_tbl2_prod_w_vector1_range7768w(0) <= vector1(20);
	wire_tbl1_tbl2_prod_w_vector1_range7779w(0) <= vector1(21);
	wire_tbl1_tbl2_prod_w_vector1_range7790w(0) <= vector1(22);
	wire_tbl1_tbl2_prod_w_vector1_range7801w(0) <= vector1(23);
	wire_tbl1_tbl2_prod_w_vector1_range7812w(0) <= vector1(24);
	wire_tbl1_tbl2_prod_w_vector1_range7823w(0) <= vector1(25);
	wire_tbl1_tbl2_prod_w_vector1_range7834w(0) <= vector1(26);
	wire_tbl1_tbl2_prod_w_vector1_range7845w(0) <= vector1(27);
	wire_tbl1_tbl2_prod_w_vector1_range7856w(0) <= vector1(28);
	wire_tbl1_tbl2_prod_w_vector1_range7867w(0) <= vector1(29);
	wire_tbl1_tbl2_prod_w_vector1_range7570w(0) <= vector1(2);
	wire_tbl1_tbl2_prod_w_vector1_range7878w(0) <= vector1(30);
	wire_tbl1_tbl2_prod_w_vector1_range7889w(0) <= vector1(31);
	wire_tbl1_tbl2_prod_w_vector1_range7900w(0) <= vector1(32);
	wire_tbl1_tbl2_prod_w_vector1_range7911w(0) <= vector1(33);
	wire_tbl1_tbl2_prod_w_vector1_range7922w(0) <= vector1(34);
	wire_tbl1_tbl2_prod_w_vector1_range7933w(0) <= vector1(35);
	wire_tbl1_tbl2_prod_w_vector1_range7944w(0) <= vector1(36);
	wire_tbl1_tbl2_prod_w_vector1_range7955w(0) <= vector1(37);
	wire_tbl1_tbl2_prod_w_vector1_range7966w(0) <= vector1(38);
	wire_tbl1_tbl2_prod_w_vector1_range7977w(0) <= vector1(39);
	wire_tbl1_tbl2_prod_w_vector1_range7581w(0) <= vector1(3);
	wire_tbl1_tbl2_prod_w_vector1_range7988w(0) <= vector1(40);
	wire_tbl1_tbl2_prod_w_vector1_range7999w(0) <= vector1(41);
	wire_tbl1_tbl2_prod_w_vector1_range8010w(0) <= vector1(42);
	wire_tbl1_tbl2_prod_w_vector1_range8021w(0) <= vector1(43);
	wire_tbl1_tbl2_prod_w_vector1_range8032w(0) <= vector1(44);
	wire_tbl1_tbl2_prod_w_vector1_range8043w(0) <= vector1(45);
	wire_tbl1_tbl2_prod_w_vector1_range8054w(0) <= vector1(46);
	wire_tbl1_tbl2_prod_w_vector1_range8065w(0) <= vector1(47);
	wire_tbl1_tbl2_prod_w_vector1_range8076w(0) <= vector1(48);
	wire_tbl1_tbl2_prod_w_vector1_range8087w(0) <= vector1(49);
	wire_tbl1_tbl2_prod_w_vector1_range7592w(0) <= vector1(4);
	wire_tbl1_tbl2_prod_w_vector1_range8098w(0) <= vector1(50);
	wire_tbl1_tbl2_prod_w_vector1_range8109w(0) <= vector1(51);
	wire_tbl1_tbl2_prod_w_vector1_range8120w(0) <= vector1(52);
	wire_tbl1_tbl2_prod_w_vector1_range8131w(0) <= vector1(53);
	wire_tbl1_tbl2_prod_w_vector1_range8142w(0) <= vector1(54);
	wire_tbl1_tbl2_prod_w_vector1_range8153w(0) <= vector1(55);
	wire_tbl1_tbl2_prod_w_vector1_range8164w(0) <= vector1(56);
	wire_tbl1_tbl2_prod_w_vector1_range8175w(0) <= vector1(57);
	wire_tbl1_tbl2_prod_w_vector1_range8186w(0) <= vector1(58);
	wire_tbl1_tbl2_prod_w_vector1_range8197w(0) <= vector1(59);
	wire_tbl1_tbl2_prod_w_vector1_range7603w(0) <= vector1(5);
	wire_tbl1_tbl2_prod_w_vector1_range8208w(0) <= vector1(60);
	wire_tbl1_tbl2_prod_w_vector1_range8219w(0) <= vector1(61);
	wire_tbl1_tbl2_prod_w_vector1_range8230w(0) <= vector1(62);
	wire_tbl1_tbl2_prod_w_vector1_range8241w(0) <= vector1(63);
	wire_tbl1_tbl2_prod_w_vector1_range8252w(0) <= vector1(64);
	wire_tbl1_tbl2_prod_w_vector1_range8263w(0) <= vector1(65);
	wire_tbl1_tbl2_prod_w_vector1_range8274w(0) <= vector1(66);
	wire_tbl1_tbl2_prod_w_vector1_range8285w(0) <= vector1(67);
	wire_tbl1_tbl2_prod_w_vector1_range8296w(0) <= vector1(68);
	wire_tbl1_tbl2_prod_w_vector1_range8307w(0) <= vector1(69);
	wire_tbl1_tbl2_prod_w_vector1_range7614w(0) <= vector1(6);
	wire_tbl1_tbl2_prod_w_vector1_range8318w(0) <= vector1(70);
	wire_tbl1_tbl2_prod_w_vector1_range8329w(0) <= vector1(71);
	wire_tbl1_tbl2_prod_w_vector1_range8340w(0) <= vector1(72);
	wire_tbl1_tbl2_prod_w_vector1_range8351w(0) <= vector1(73);
	wire_tbl1_tbl2_prod_w_vector1_range8362w(0) <= vector1(74);
	wire_tbl1_tbl2_prod_w_vector1_range8373w(0) <= vector1(75);
	wire_tbl1_tbl2_prod_w_vector1_range8384w(0) <= vector1(76);
	wire_tbl1_tbl2_prod_w_vector1_range8395w(0) <= vector1(77);
	wire_tbl1_tbl2_prod_w_vector1_range8406w(0) <= vector1(78);
	wire_tbl1_tbl2_prod_w_vector1_range8417w(0) <= vector1(79);
	wire_tbl1_tbl2_prod_w_vector1_range7625w(0) <= vector1(7);
	wire_tbl1_tbl2_prod_w_vector1_range8428w(0) <= vector1(80);
	wire_tbl1_tbl2_prod_w_vector1_range8439w(0) <= vector1(81);
	wire_tbl1_tbl2_prod_w_vector1_range8450w(0) <= vector1(82);
	wire_tbl1_tbl2_prod_w_vector1_range8461w(0) <= vector1(83);
	wire_tbl1_tbl2_prod_w_vector1_range8472w(0) <= vector1(84);
	wire_tbl1_tbl2_prod_w_vector1_range8483w(0) <= vector1(85);
	wire_tbl1_tbl2_prod_w_vector1_range8494w(0) <= vector1(86);
	wire_tbl1_tbl2_prod_w_vector1_range8505w(0) <= vector1(87);
	wire_tbl1_tbl2_prod_w_vector1_range8516w(0) <= vector1(88);
	wire_tbl1_tbl2_prod_w_vector1_range8527w(0) <= vector1(89);
	wire_tbl1_tbl2_prod_w_vector1_range7636w(0) <= vector1(8);
	wire_tbl1_tbl2_prod_w_vector1_range8538w(0) <= vector1(90);
	wire_tbl1_tbl2_prod_w_vector1_range8549w(0) <= vector1(91);
	wire_tbl1_tbl2_prod_w_vector1_range7647w(0) <= vector1(9);
	wire_tbl1_tbl2_prod_w_vector2_range6619w(0) <= vector2(0);
	wire_tbl1_tbl2_prod_w_vector2_range6721w(0) <= vector2(10);
	wire_tbl1_tbl2_prod_w_vector2_range6731w(0) <= vector2(11);
	wire_tbl1_tbl2_prod_w_vector2_range6741w(0) <= vector2(12);
	wire_tbl1_tbl2_prod_w_vector2_range6751w(0) <= vector2(13);
	wire_tbl1_tbl2_prod_w_vector2_range6761w(0) <= vector2(14);
	wire_tbl1_tbl2_prod_w_vector2_range6771w(0) <= vector2(15);
	wire_tbl1_tbl2_prod_w_vector2_range6781w(0) <= vector2(16);
	wire_tbl1_tbl2_prod_w_vector2_range6791w(0) <= vector2(17);
	wire_tbl1_tbl2_prod_w_vector2_range6801w(0) <= vector2(18);
	wire_tbl1_tbl2_prod_w_vector2_range6811w(0) <= vector2(19);
	wire_tbl1_tbl2_prod_w_vector2_range6631w(0) <= vector2(1);
	wire_tbl1_tbl2_prod_w_vector2_range6821w(0) <= vector2(20);
	wire_tbl1_tbl2_prod_w_vector2_range6831w(0) <= vector2(21);
	wire_tbl1_tbl2_prod_w_vector2_range6841w(0) <= vector2(22);
	wire_tbl1_tbl2_prod_w_vector2_range6851w(0) <= vector2(23);
	wire_tbl1_tbl2_prod_w_vector2_range6861w(0) <= vector2(24);
	wire_tbl1_tbl2_prod_w_vector2_range6871w(0) <= vector2(25);
	wire_tbl1_tbl2_prod_w_vector2_range6881w(0) <= vector2(26);
	wire_tbl1_tbl2_prod_w_vector2_range6891w(0) <= vector2(27);
	wire_tbl1_tbl2_prod_w_vector2_range6901w(0) <= vector2(28);
	wire_tbl1_tbl2_prod_w_vector2_range6911w(0) <= vector2(29);
	wire_tbl1_tbl2_prod_w_vector2_range6641w(0) <= vector2(2);
	wire_tbl1_tbl2_prod_w_vector2_range6921w(0) <= vector2(30);
	wire_tbl1_tbl2_prod_w_vector2_range6931w(0) <= vector2(31);
	wire_tbl1_tbl2_prod_w_vector2_range6941w(0) <= vector2(32);
	wire_tbl1_tbl2_prod_w_vector2_range6951w(0) <= vector2(33);
	wire_tbl1_tbl2_prod_w_vector2_range6961w(0) <= vector2(34);
	wire_tbl1_tbl2_prod_w_vector2_range6971w(0) <= vector2(35);
	wire_tbl1_tbl2_prod_w_vector2_range6981w(0) <= vector2(36);
	wire_tbl1_tbl2_prod_w_vector2_range6991w(0) <= vector2(37);
	wire_tbl1_tbl2_prod_w_vector2_range7001w(0) <= vector2(38);
	wire_tbl1_tbl2_prod_w_vector2_range7011w(0) <= vector2(39);
	wire_tbl1_tbl2_prod_w_vector2_range6651w(0) <= vector2(3);
	wire_tbl1_tbl2_prod_w_vector2_range7021w(0) <= vector2(40);
	wire_tbl1_tbl2_prod_w_vector2_range7031w(0) <= vector2(41);
	wire_tbl1_tbl2_prod_w_vector2_range7041w(0) <= vector2(42);
	wire_tbl1_tbl2_prod_w_vector2_range7051w(0) <= vector2(43);
	wire_tbl1_tbl2_prod_w_vector2_range7061w(0) <= vector2(44);
	wire_tbl1_tbl2_prod_w_vector2_range7071w(0) <= vector2(45);
	wire_tbl1_tbl2_prod_w_vector2_range7081w(0) <= vector2(46);
	wire_tbl1_tbl2_prod_w_vector2_range7091w(0) <= vector2(47);
	wire_tbl1_tbl2_prod_w_vector2_range7101w(0) <= vector2(48);
	wire_tbl1_tbl2_prod_w_vector2_range7111w(0) <= vector2(49);
	wire_tbl1_tbl2_prod_w_vector2_range6661w(0) <= vector2(4);
	wire_tbl1_tbl2_prod_w_vector2_range7121w(0) <= vector2(50);
	wire_tbl1_tbl2_prod_w_vector2_range7131w(0) <= vector2(51);
	wire_tbl1_tbl2_prod_w_vector2_range7141w(0) <= vector2(52);
	wire_tbl1_tbl2_prod_w_vector2_range7151w(0) <= vector2(53);
	wire_tbl1_tbl2_prod_w_vector2_range7161w(0) <= vector2(54);
	wire_tbl1_tbl2_prod_w_vector2_range7171w(0) <= vector2(55);
	wire_tbl1_tbl2_prod_w_vector2_range7181w(0) <= vector2(56);
	wire_tbl1_tbl2_prod_w_vector2_range7191w(0) <= vector2(57);
	wire_tbl1_tbl2_prod_w_vector2_range7201w(0) <= vector2(58);
	wire_tbl1_tbl2_prod_w_vector2_range7211w(0) <= vector2(59);
	wire_tbl1_tbl2_prod_w_vector2_range6671w(0) <= vector2(5);
	wire_tbl1_tbl2_prod_w_vector2_range7221w(0) <= vector2(60);
	wire_tbl1_tbl2_prod_w_vector2_range7231w(0) <= vector2(61);
	wire_tbl1_tbl2_prod_w_vector2_range7241w(0) <= vector2(62);
	wire_tbl1_tbl2_prod_w_vector2_range7251w(0) <= vector2(63);
	wire_tbl1_tbl2_prod_w_vector2_range7261w(0) <= vector2(64);
	wire_tbl1_tbl2_prod_w_vector2_range7271w(0) <= vector2(65);
	wire_tbl1_tbl2_prod_w_vector2_range7281w(0) <= vector2(66);
	wire_tbl1_tbl2_prod_w_vector2_range7291w(0) <= vector2(67);
	wire_tbl1_tbl2_prod_w_vector2_range7301w(0) <= vector2(68);
	wire_tbl1_tbl2_prod_w_vector2_range7311w(0) <= vector2(69);
	wire_tbl1_tbl2_prod_w_vector2_range6681w(0) <= vector2(6);
	wire_tbl1_tbl2_prod_w_vector2_range7321w(0) <= vector2(70);
	wire_tbl1_tbl2_prod_w_vector2_range7331w(0) <= vector2(71);
	wire_tbl1_tbl2_prod_w_vector2_range7341w(0) <= vector2(72);
	wire_tbl1_tbl2_prod_w_vector2_range7351w(0) <= vector2(73);
	wire_tbl1_tbl2_prod_w_vector2_range7361w(0) <= vector2(74);
	wire_tbl1_tbl2_prod_w_vector2_range7371w(0) <= vector2(75);
	wire_tbl1_tbl2_prod_w_vector2_range7381w(0) <= vector2(76);
	wire_tbl1_tbl2_prod_w_vector2_range7391w(0) <= vector2(77);
	wire_tbl1_tbl2_prod_w_vector2_range7401w(0) <= vector2(78);
	wire_tbl1_tbl2_prod_w_vector2_range7411w(0) <= vector2(79);
	wire_tbl1_tbl2_prod_w_vector2_range6691w(0) <= vector2(7);
	wire_tbl1_tbl2_prod_w_vector2_range7421w(0) <= vector2(80);
	wire_tbl1_tbl2_prod_w_vector2_range7431w(0) <= vector2(81);
	wire_tbl1_tbl2_prod_w_vector2_range7441w(0) <= vector2(82);
	wire_tbl1_tbl2_prod_w_vector2_range7451w(0) <= vector2(83);
	wire_tbl1_tbl2_prod_w_vector2_range7461w(0) <= vector2(84);
	wire_tbl1_tbl2_prod_w_vector2_range7471w(0) <= vector2(85);
	wire_tbl1_tbl2_prod_w_vector2_range7481w(0) <= vector2(86);
	wire_tbl1_tbl2_prod_w_vector2_range7491w(0) <= vector2(87);
	wire_tbl1_tbl2_prod_w_vector2_range7501w(0) <= vector2(88);
	wire_tbl1_tbl2_prod_w_vector2_range7511w(0) <= vector2(89);
	wire_tbl1_tbl2_prod_w_vector2_range6701w(0) <= vector2(8);
	wire_tbl1_tbl2_prod_w_vector2_range7521w(0) <= vector2(90);
	wire_tbl1_tbl2_prod_w_vector2_range7531w(0) <= vector2(91);
	wire_tbl1_tbl2_prod_w_vector2_range6711w(0) <= vector2(9);
	sum :  ALTFP_EXa_altmult_opt_csa_nsf
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => car_two_wo,
		datab => sum_two_wo,
		result => wire_sum_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN car_two_adj_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN car_two_adj_reg0 <= car_two_adj;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg0 <= lowest_bits_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg1 <= lowest_bits_wi_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg2 <= lowest_bits_wi_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lsb_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lsb_prod_wi_reg0 <= lsb_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mid_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mid_prod_wi_reg0 <= mid_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN msb_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN msb_prod_wi_reg0 <= msb_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sum_two_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sum_two_reg0 <= sum_two;
			END IF;
		END IF;
	END PROCESS;
	wire_compress_a_dataa <= ( "0" & wire_a(60 DOWNTO 31));
	compress_a :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		cout => wire_compress_a_cout,
		dataa => wire_compress_a_dataa,
		datab => wire_a(30 DOWNTO 0),
		result => wire_compress_a_result
	  );
	wire_compress_b_dataa <= ( "0" & wire_b(60 DOWNTO 31));
	compress_b :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		cout => wire_compress_b_cout,
		dataa => wire_compress_b_dataa,
		datab => wire_b(30 DOWNTO 0),
		result => wire_compress_b_result
	  );
	lsb_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 31,
		LPM_WIDTHB => 31,
		LPM_WIDTHP => 62,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_a(30 DOWNTO 0),
		datab => wire_b(30 DOWNTO 0),
		result => wire_lsb_prod_result
	  );
	wire_mid_prod_dataa <= ( wire_compress_a_cout & wire_compress_a_result);
	wire_mid_prod_datab <= ( wire_compress_b_cout & wire_compress_b_result);
	mid_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 32,
		LPM_WIDTHB => 32,
		LPM_WIDTHP => 64,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_mid_prod_dataa,
		datab => wire_mid_prod_datab,
		result => wire_mid_prod_result
	  );
	wire_msb_prod_dataa <= ( "0" & wire_a(60 DOWNTO 31));
	msb_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 31,
		LPM_WIDTHB => 30,
		LPM_WIDTHP => 61,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_msb_prod_dataa,
		datab => wire_b(60 DOWNTO 31),
		result => wire_msb_prod_result
	  );

 END RTL; --ALTFP_EXa_altmult_opt_45e


--altmult_opt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" LPM_PIPELINE=5 LPM_WIDTHA=61 LPM_WIDTHB=59 LPM_WIDTHP=120 aclr clken clock dataa datab result
--VERSION_BEGIN 16.0 cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END


--altmult_opt_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=2 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=90 aclr clken clock dataa datab result
--VERSION_BEGIN 16.0 cbx_altmult_opt 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_mult 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_padd 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altmult_opt_csa_lsf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (89 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (89 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (89 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altmult_opt_csa_lsf;

 ARCHITECTURE RTL OF ALTFP_EXa_altmult_opt_csa_lsf IS

	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub3_result;
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 90
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub3_result
	  );

 END RTL; --ALTFP_EXa_altmult_opt_csa_lsf

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 lpm_mult 3 reg 458 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altmult_opt_95e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (60 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (58 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (119 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altmult_opt_95e;

 ARCHITECTURE RTL OF ALTFP_EXa_altmult_opt_95e IS

	 SIGNAL  wire_sum_result	:	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL	 car_two_adj_reg0	:	STD_LOGIC_VECTOR(89 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg0	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg1	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_bits_wi_reg2	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lsb_prod_wi_reg0	:	STD_LOGIC_VECTOR(61 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mid_prod_wi_reg0	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 msb_prod_wi_reg0	:	STD_LOGIC_VECTOR(58 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sum_two_reg0	:	STD_LOGIC_VECTOR(89 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_compress_a_cout	:	STD_LOGIC;
	 SIGNAL  wire_compress_a_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_compress_a_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_compress_b_cout	:	STD_LOGIC;
	 SIGNAL  wire_compress_b_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_compress_b_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_lsb_prod_result	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_mid_prod_dataa	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_mid_prod_datab	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_mid_prod_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_msb_prod_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_msb_prod_result	:	STD_LOGIC_VECTOR (58 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9079w9088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9019w9189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9013w9199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9007w9209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9001w9219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8995w9229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8989w9239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8983w9249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8977w9259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8971w9269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8965w9279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9073w9099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8959w9289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8953w9299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8947w9309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8941w9319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8935w9329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8929w9339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8923w9349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8917w9359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8911w9369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8905w9379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9067w9109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8899w9389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8893w9399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8887w9409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8881w9419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8875w9429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8869w9439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8863w9449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8857w9459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8851w9469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8845w9479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9061w9119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8839w9489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8833w9499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8827w9509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8821w9519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8815w9529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8809w9539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8803w9549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8797w9559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8791w9569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8785w9579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9055w9129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8779w9589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8773w9599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8767w9609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8761w9619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8755w9629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8749w9639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8743w9649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8737w9659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8731w9669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8724w9679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9049w9139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8719w9689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8714w9699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8710w9709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8706w9719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8702w9729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8698w9739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8694w9749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8690w9759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8686w9769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8682w9779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9043w9149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8678w9789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8674w9799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8670w9809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8666w9819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8662w9829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8658w9839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8654w9849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8650w9859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8646w9869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8642w9879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9037w9159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8638w9889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8634w9899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8630w9909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8626w9919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8622w9929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8618w9939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8614w9949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8610w9959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8606w9969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8600w9979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9031w9169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9025w9179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9086w9995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9188w10106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9198w10117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9208w10128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9218w10139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9228w10150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9238w10161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9248w10172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9258w10183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9268w10194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9278w10205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9098w10007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9288w10216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9298w10227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9308w10238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9318w10249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9328w10260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9338w10271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9348w10282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9358w10293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9368w10304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9378w10315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9108w10018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9388w10326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9398w10337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9408w10348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9418w10359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9428w10370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9438w10381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9448w10392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9458w10403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9468w10414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9478w10425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9118w10029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9488w10436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9498w10447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9508w10458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9518w10469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9528w10480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9538w10491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9548w10502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9558w10513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9568w10524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9578w10535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9128w10040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9588w10546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9598w10557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9608w10568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9618w10579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9628w10590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9638w10601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9648w10612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9658w10623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9668w10634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9678w10645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9138w10051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9688w10656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9698w10667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9708w10678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9718w10689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9728w10700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9738w10711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9748w10722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9758w10733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9768w10744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9778w10755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9148w10062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9788w10766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9798w10777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9808w10788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9818w10799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9828w10810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9838w10821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9848w10832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9858w10843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9868w10854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9878w10865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9158w10073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9888w10876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9898w10887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9908w10898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9918w10909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9928w10920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9938w10931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9948w10942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9958w10953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9968w10964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9978w10975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9168w10084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_sum_one_range9178w10095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9080w9081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9020w9021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9014w9015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9008w9009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9002w9003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8996w8997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8990w8991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8984w8985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8978w8979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8972w8973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8966w8967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9074w9075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8960w8961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8954w8955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8948w8949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8942w8943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8936w8937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8930w8931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8924w8925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8918w8919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8912w8913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8906w8907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9068w9069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8900w8901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8894w8895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8888w8889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8882w8883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8876w8877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8870w8871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8864w8865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8858w8859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8852w8853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8846w8847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9062w9063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8840w8841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8834w8835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8828w8829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8822w8823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8816w8817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8810w8811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8804w8805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8798w8799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8792w8793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8786w8787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9056w9057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8780w8781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8774w8775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8768w8769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8762w8763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8756w8757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8750w8751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8744w8745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8738w8739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8732w8733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8726w8727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9050w9051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8721w8722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8716w8717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9044w9045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9038w9039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9032w9033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9026w9027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9077w9078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9017w9018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9011w9012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9005w9006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8999w9000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8993w8994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8987w8988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8981w8982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8975w8976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8969w8970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8963w8964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9071w9072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8957w8958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8951w8952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8945w8946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8939w8940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8933w8934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8927w8928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8921w8922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8915w8916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8909w8910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8903w8904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9065w9066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8897w8898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8891w8892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8885w8886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8879w8880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8873w8874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8867w8868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8861w8862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8855w8856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8849w8850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8843w8844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9059w9060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8837w8838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8831w8832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8825w8826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8819w8820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8813w8814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8807w8808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8801w8802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8795w8796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8789w8790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8783w8784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9053w9054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8777w8778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8771w8772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8765w8766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8759w8760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8753w8754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8747w8748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8741w8742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8735w8736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8729w8730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9047w9048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9041w9042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9035w9036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9029w9030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9023w9024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range9990w9997w9998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10102w10108w10109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10113w10119w10120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10124w10130w10131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10135w10141w10142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10146w10152w10153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10157w10163w10164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10168w10174w10175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10179w10185w10186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10190w10196w10197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10201w10207w10208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10003w10009w10010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10212w10218w10219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10223w10229w10230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10234w10240w10241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10245w10251w10252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10256w10262w10263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10267w10273w10274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10278w10284w10285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10289w10295w10296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10300w10306w10307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10311w10317w10318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10014w10020w10021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10322w10328w10329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10333w10339w10340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10344w10350w10351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10355w10361w10362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10366w10372w10373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10377w10383w10384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10388w10394w10395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10399w10405w10406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10410w10416w10417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10421w10427w10428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10025w10031w10032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10432w10438w10439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10443w10449w10450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10454w10460w10461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10465w10471w10472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10476w10482w10483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10487w10493w10494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10498w10504w10505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10509w10515w10516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10520w10526w10527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10531w10537w10538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10036w10042w10043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10542w10548w10549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10553w10559w10560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10564w10570w10571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10575w10581w10582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10586w10592w10593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10597w10603w10604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10608w10614w10615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10619w10625w10626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10630w10636w10637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10641w10647w10648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10047w10053w10054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10652w10658w10659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10663w10669w10670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10674w10680w10681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10685w10691w10692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10696w10702w10703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10707w10713w10714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10718w10724w10725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10729w10735w10736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10740w10746w10747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10751w10757w10758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10058w10064w10065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10762w10768w10769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10773w10779w10780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10784w10790w10791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10795w10801w10802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10806w10812w10813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10817w10823w10824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10828w10834w10835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10839w10845w10846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10850w10856w10857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10861w10867w10868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10069w10075w10076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10872w10878w10879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10883w10889w10890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10894w10900w10901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10905w10911w10912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10916w10922w10923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10927w10933w10934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10938w10944w10945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10949w10955w10956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10960w10966w10967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10971w10977w10978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10080w10086w10087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10091w10097w10098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9083w9090w9091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9185w9191w9192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9195w9201w9202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9205w9211w9212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9215w9221w9222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9225w9231w9232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9235w9241w9242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9245w9251w9252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9255w9261w9262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9265w9271w9272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9275w9281w9282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9095w9101w9102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9285w9291w9292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9295w9301w9302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9305w9311w9312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9315w9321w9322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9325w9331w9332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9335w9341w9342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9345w9351w9352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9355w9361w9362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9365w9371w9372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9375w9381w9382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9105w9111w9112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9385w9391w9392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9395w9401w9402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9405w9411w9412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9415w9421w9422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9425w9431w9432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9435w9441w9442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9445w9451w9452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9455w9461w9462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9465w9471w9472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9475w9481w9482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9115w9121w9122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9485w9491w9492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9495w9501w9502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9505w9511w9512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9515w9521w9522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9525w9531w9532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9535w9541w9542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9545w9551w9552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9555w9561w9562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9565w9571w9572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9575w9581w9582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9125w9131w9132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9585w9591w9592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9595w9601w9602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9605w9611w9612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9615w9621w9622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9625w9631w9632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9635w9641w9642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9645w9651w9652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9655w9661w9662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9665w9671w9672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9675w9681w9682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9135w9141w9142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9685w9691w9692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9695w9701w9702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9705w9711w9712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9715w9721w9722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9725w9731w9732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9735w9741w9742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9745w9751w9752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9755w9761w9762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9765w9771w9772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9775w9781w9782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9145w9151w9152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9785w9791w9792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9795w9801w9802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9805w9811w9812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9815w9821w9822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9825w9831w9832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9835w9841w9842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9845w9851w9852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9855w9861w9862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9865w9871w9872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9875w9881w9882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9155w9161w9162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9885w9891w9892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9895w9901w9902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9905w9911w9912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9915w9921w9922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9925w9931w9932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9935w9941w9942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9945w9951w9952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9955w9961w9962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9965w9971w9972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9975w9981w9982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9165w9171w9172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9175w9181w9182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector1_range9990w9997w9998w9999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w10099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9083w9090w9091w9092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9185w9191w9192w9193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9195w9201w9202w9203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9205w9211w9212w9213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9215w9221w9222w9223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9225w9231w9232w9233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9235w9241w9242w9243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9245w9251w9252w9253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9255w9261w9262w9263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9265w9271w9272w9273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9275w9281w9282w9283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9095w9101w9102w9103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9285w9291w9292w9293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9295w9301w9302w9303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9305w9311w9312w9313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9315w9321w9322w9323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9325w9331w9332w9333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9335w9341w9342w9343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9345w9351w9352w9353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9355w9361w9362w9363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9365w9371w9372w9373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9375w9381w9382w9383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9105w9111w9112w9113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9385w9391w9392w9393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9395w9401w9402w9403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9405w9411w9412w9413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9415w9421w9422w9423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9425w9431w9432w9433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9435w9441w9442w9443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9445w9451w9452w9453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9455w9461w9462w9463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9465w9471w9472w9473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9475w9481w9482w9483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9115w9121w9122w9123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9485w9491w9492w9493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9495w9501w9502w9503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9505w9511w9512w9513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9515w9521w9522w9523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9525w9531w9532w9533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9535w9541w9542w9543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9545w9551w9552w9553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9555w9561w9562w9563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9565w9571w9572w9573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9575w9581w9582w9583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9125w9131w9132w9133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9585w9591w9592w9593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9595w9601w9602w9603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9605w9611w9612w9613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9615w9621w9622w9623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9625w9631w9632w9633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9635w9641w9642w9643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9645w9651w9652w9653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9655w9661w9662w9663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9665w9671w9672w9673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9675w9681w9682w9683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9135w9141w9142w9143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9685w9691w9692w9693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9695w9701w9702w9703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9705w9711w9712w9713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9715w9721w9722w9723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9725w9731w9732w9733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9735w9741w9742w9743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9745w9751w9752w9753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9755w9761w9762w9763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9765w9771w9772w9773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9775w9781w9782w9783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9145w9151w9152w9153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9785w9791w9792w9793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9795w9801w9802w9803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9805w9811w9812w9813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9815w9821w9822w9823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9825w9831w9832w9833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9835w9841w9842w9843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9845w9851w9852w9853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9855w9861w9862w9863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9865w9871w9872w9873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9875w9881w9882w9883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9155w9161w9162w9163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9885w9891w9892w9893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9895w9901w9902w9903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9905w9911w9912w9913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9915w9921w9922w9923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9925w9931w9932w9933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9935w9941w9942w9943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9945w9951w9952w9953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9955w9961w9962w9963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9965w9971w9972w9973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9975w9981w9982w9983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9165w9171w9172w9173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9175w9181w9182w9183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range9990w9991w9992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10102w10103w10104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10113w10114w10115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10124w10125w10126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10135w10136w10137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10146w10147w10148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10157w10158w10159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10168w10169w10170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10179w10180w10181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10190w10191w10192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10201w10202w10203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10003w10004w10005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10212w10213w10214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10223w10224w10225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10234w10235w10236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10245w10246w10247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10256w10257w10258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10267w10268w10269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10278w10279w10280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10289w10290w10291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10300w10301w10302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10311w10312w10313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10014w10015w10016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10322w10323w10324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10333w10334w10335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10344w10345w10346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10355w10356w10357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10366w10367w10368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10377w10378w10379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10388w10389w10390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10399w10400w10401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10410w10411w10412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10421w10422w10423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10025w10026w10027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10432w10433w10434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10443w10444w10445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10454w10455w10456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10465w10466w10467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10476w10477w10478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10487w10488w10489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10498w10499w10500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10509w10510w10511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10520w10521w10522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10531w10532w10533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10036w10037w10038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10542w10543w10544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10553w10554w10555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10564w10565w10566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10575w10576w10577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10586w10587w10588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10597w10598w10599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10608w10609w10610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10619w10620w10621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10630w10631w10632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10641w10642w10643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10047w10048w10049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10652w10653w10654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10663w10664w10665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10674w10675w10676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10685w10686w10687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10696w10697w10698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10707w10708w10709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10718w10719w10720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10729w10730w10731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10740w10741w10742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10751w10752w10753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10058w10059w10060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10762w10763w10764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10773w10774w10775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10784w10785w10786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10795w10796w10797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10806w10807w10808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10817w10818w10819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10828w10829w10830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10839w10840w10841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10850w10851w10852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10861w10862w10863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10069w10070w10071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10872w10873w10874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10883w10884w10885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10894w10895w10896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10905w10906w10907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10916w10917w10918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10927w10928w10929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10938w10939w10940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10949w10950w10951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10960w10961w10962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10971w10972w10973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10080w10081w10082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10091w10092w10093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9083w9084w9085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9185w9186w9187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9195w9196w9197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9205w9206w9207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9215w9216w9217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9225w9226w9227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9235w9236w9237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9245w9246w9247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9255w9256w9257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9265w9266w9267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9275w9276w9277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9095w9096w9097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9285w9286w9287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9295w9296w9297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9305w9306w9307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9315w9316w9317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9325w9326w9327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9335w9336w9337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9345w9346w9347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9355w9356w9357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9365w9366w9367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9375w9376w9377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9105w9106w9107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9385w9386w9387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9395w9396w9397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9405w9406w9407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9415w9416w9417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9425w9426w9427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9435w9436w9437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9445w9446w9447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9455w9456w9457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9465w9466w9467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9475w9476w9477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9115w9116w9117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9485w9486w9487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9495w9496w9497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9505w9506w9507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9515w9516w9517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9525w9526w9527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9535w9536w9537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9545w9546w9547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9555w9556w9557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9565w9566w9567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9575w9576w9577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9125w9126w9127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9585w9586w9587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9595w9596w9597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9605w9606w9607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9615w9616w9617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9625w9626w9627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9635w9636w9637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9645w9646w9647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9655w9656w9657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9665w9666w9667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9675w9676w9677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9135w9136w9137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9685w9686w9687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9695w9696w9697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9705w9706w9707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9715w9716w9717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9725w9726w9727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9735w9736w9737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9745w9746w9747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9755w9756w9757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9765w9766w9767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9775w9776w9777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9145w9146w9147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9785w9786w9787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9795w9796w9797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9805w9806w9807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9815w9816w9817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9825w9826w9827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9835w9836w9837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9845w9846w9847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9855w9856w9857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9865w9866w9867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9875w9876w9877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9155w9156w9157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9885w9886w9887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9895w9896w9897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9905w9906w9907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9915w9916w9917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9925w9926w9927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9935w9936w9937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9945w9946w9947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9955w9956w9957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9965w9966w9967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9975w9976w9977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9165w9166w9167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9175w9176w9177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  car_one :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_one_adj :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_two :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_two_adj :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  car_two_wo :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  lowest_bits_wi :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lowest_bits_wo :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lsb_prod_wi :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  lsb_prod_wo :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  mid_prod_wi :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  mid_prod_wo :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  msb_prod_out :	STD_LOGIC_VECTOR (58 DOWNTO 0);
	 SIGNAL  msb_prod_wi :	STD_LOGIC_VECTOR (58 DOWNTO 0);
	 SIGNAL  msb_prod_wo :	STD_LOGIC_VECTOR (58 DOWNTO 0);
	 SIGNAL  neg_lsb :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  neg_msb :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  sum_one :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  sum_two :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  sum_two_wo :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  vector1 :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  vector2 :	STD_LOGIC_VECTOR (89 DOWNTO 0);
	 SIGNAL  wire_a :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  wire_b :	STD_LOGIC_VECTOR (58 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range9988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_car_one_adj_range10090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range8716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_lsb_prod_wo_range9026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range8729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_msb_prod_wo_range9023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range8603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_lsb_range9028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range8600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_neg_msb_range9025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_sum_one_range9178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range9990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector1_range10091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_w_vector2_range9175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  ALTFP_EXa_altmult_opt_csa_lsf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(89 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(89 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(89 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9079w9088w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9079w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9082w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9019w9189w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9019w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9022w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9013w9199w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9013w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9016w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9007w9209w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9007w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9010w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9001w9219w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9001w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9004w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8995w9229w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8995w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8998w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8989w9239w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8989w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8992w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8983w9249w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8983w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8986w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8977w9259w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8977w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8980w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8971w9269w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8971w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8974w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8965w9279w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8965w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8968w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9073w9099w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9073w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9076w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8959w9289w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8959w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8962w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8953w9299w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8953w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8956w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8947w9309w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8947w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8950w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8941w9319w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8941w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8944w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8935w9329w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8935w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8938w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8929w9339w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8929w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8932w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8923w9349w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8923w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8926w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8917w9359w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8917w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8920w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8911w9369w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8911w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8914w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8905w9379w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8905w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8908w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9067w9109w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9067w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9070w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8899w9389w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8899w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8902w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8893w9399w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8893w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8896w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8887w9409w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8887w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8890w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8881w9419w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8881w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8884w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8875w9429w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8875w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8878w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8869w9439w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8869w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8872w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8863w9449w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8863w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8866w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8857w9459w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8857w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8860w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8851w9469w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8851w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8854w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8845w9479w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8845w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8848w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9061w9119w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9061w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9064w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8839w9489w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8839w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8842w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8833w9499w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8833w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8836w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8827w9509w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8827w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8830w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8821w9519w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8821w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8824w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8815w9529w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8815w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8818w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8809w9539w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8809w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8812w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8803w9549w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8803w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8806w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8797w9559w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8797w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8800w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8791w9569w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8791w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8794w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8785w9579w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8785w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8788w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9055w9129w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9055w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9058w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8779w9589w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8779w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8782w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8773w9599w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8773w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8776w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8767w9609w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8767w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8770w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8761w9619w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8761w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8764w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8755w9629w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8755w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8758w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8749w9639w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8749w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8752w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8743w9649w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8743w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8746w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8737w9659w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8737w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8740w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8731w9669w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8731w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8734w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8724w9679w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8724w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8728w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9049w9139w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9049w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9052w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8719w9689w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8719w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8723w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8714w9699w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8714w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8718w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8710w9709w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8710w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8712w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8706w9719w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8706w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8708w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8702w9729w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8702w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8704w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8698w9739w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8698w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8700w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8694w9749w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8694w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8696w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8690w9759w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8690w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8692w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8686w9769w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8686w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8688w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8682w9779w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8682w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8684w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9043w9149w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9043w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9046w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8678w9789w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8678w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8680w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8674w9799w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8674w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8676w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8670w9809w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8670w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8672w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8666w9819w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8666w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8668w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8662w9829w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8662w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8664w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8658w9839w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8658w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8660w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8654w9849w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8654w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8656w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8650w9859w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8650w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8652w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8646w9869w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8646w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8648w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8642w9879w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8642w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8644w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9037w9159w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9037w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9040w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8638w9889w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8638w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8640w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8634w9899w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8634w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8636w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8630w9909w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8630w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8632w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8626w9919w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8626w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8628w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8622w9929w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8622w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8624w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8618w9939w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8618w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8620w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8614w9949w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8614w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8616w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8610w9959w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8610w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8612w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8606w9969w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8606w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8608w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8600w9979w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range8600w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8603w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9031w9169w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9031w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9034w(0);
	wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9025w9179w(0) <= wire_tbl3_taylor_prod_w_neg_msb_range9025w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9028w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9086w9995w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9086w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range9988w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9188w10106w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9188w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10101w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9198w10117w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9198w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10112w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9208w10128w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9208w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10123w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9218w10139w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9218w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10134w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9228w10150w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9228w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10145w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9238w10161w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9238w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10156w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9248w10172w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9248w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10167w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9258w10183w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9258w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10178w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9268w10194w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9268w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10189w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9278w10205w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9278w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10200w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9098w10007w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9098w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10002w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9288w10216w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9288w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10211w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9298w10227w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9298w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10222w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9308w10238w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9308w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10233w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9318w10249w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9318w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10244w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9328w10260w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9328w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10255w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9338w10271w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9338w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10266w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9348w10282w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9348w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10277w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9358w10293w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9358w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10288w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9368w10304w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9368w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10299w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9378w10315w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9378w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10310w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9108w10018w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9108w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10013w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9388w10326w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9388w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10321w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9398w10337w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9398w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10332w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9408w10348w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9408w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10343w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9418w10359w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9418w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10354w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9428w10370w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9428w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10365w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9438w10381w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9438w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10376w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9448w10392w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9448w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10387w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9458w10403w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9458w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10398w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9468w10414w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9468w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10409w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9478w10425w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9478w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10420w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9118w10029w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9118w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10024w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9488w10436w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9488w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10431w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9498w10447w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9498w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10442w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9508w10458w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9508w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10453w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9518w10469w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9518w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10464w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9528w10480w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9528w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10475w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9538w10491w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9538w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10486w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9548w10502w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9548w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10497w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9558w10513w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9558w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10508w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9568w10524w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9568w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10519w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9578w10535w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9578w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10530w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9128w10040w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9128w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10035w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9588w10546w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9588w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10541w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9598w10557w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9598w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10552w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9608w10568w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9608w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10563w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9618w10579w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9618w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10574w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9628w10590w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9628w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10585w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9638w10601w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9638w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10596w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9648w10612w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9648w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10607w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9658w10623w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9658w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10618w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9668w10634w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9668w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10629w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9678w10645w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9678w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10640w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9138w10051w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9138w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10046w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9688w10656w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9688w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10651w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9698w10667w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9698w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10662w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9708w10678w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9708w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10673w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9718w10689w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9718w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10684w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9728w10700w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9728w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10695w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9738w10711w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9738w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10706w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9748w10722w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9748w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10717w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9758w10733w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9758w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10728w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9768w10744w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9768w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10739w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9778w10755w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9778w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10750w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9148w10062w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9148w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10057w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9788w10766w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9788w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10761w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9798w10777w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9798w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10772w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9808w10788w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9808w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10783w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9818w10799w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9818w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10794w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9828w10810w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9828w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10805w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9838w10821w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9838w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10816w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9848w10832w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9848w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10827w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9858w10843w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9858w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10838w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9868w10854w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9868w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10849w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9878w10865w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9878w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10860w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9158w10073w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9158w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10068w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9888w10876w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9888w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10871w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9898w10887w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9898w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10882w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9908w10898w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9908w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10893w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9918w10909w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9918w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10904w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9928w10920w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9928w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10915w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9938w10931w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9938w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10926w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9948w10942w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9948w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10937w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9958w10953w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9958w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10948w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9968w10964w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9968w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10959w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9978w10975w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9978w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10970w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9168w10084w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9168w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10079w(0);
	wire_tbl3_taylor_prod_w_lg_w_sum_one_range9178w10095w(0) <= wire_tbl3_taylor_prod_w_sum_one_range9178w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10090w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9996w(0) <= wire_tbl3_taylor_prod_w_vector1_range9990w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range9988w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9997w(0) <= wire_tbl3_taylor_prod_w_vector1_range9990w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9086w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10107w(0) <= wire_tbl3_taylor_prod_w_vector1_range10102w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10101w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10108w(0) <= wire_tbl3_taylor_prod_w_vector1_range10102w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9188w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10118w(0) <= wire_tbl3_taylor_prod_w_vector1_range10113w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10112w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10119w(0) <= wire_tbl3_taylor_prod_w_vector1_range10113w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9198w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10129w(0) <= wire_tbl3_taylor_prod_w_vector1_range10124w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10123w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10130w(0) <= wire_tbl3_taylor_prod_w_vector1_range10124w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9208w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10140w(0) <= wire_tbl3_taylor_prod_w_vector1_range10135w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10134w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10141w(0) <= wire_tbl3_taylor_prod_w_vector1_range10135w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9218w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10151w(0) <= wire_tbl3_taylor_prod_w_vector1_range10146w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10145w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10152w(0) <= wire_tbl3_taylor_prod_w_vector1_range10146w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9228w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10162w(0) <= wire_tbl3_taylor_prod_w_vector1_range10157w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10156w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10163w(0) <= wire_tbl3_taylor_prod_w_vector1_range10157w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9238w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10173w(0) <= wire_tbl3_taylor_prod_w_vector1_range10168w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10167w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10174w(0) <= wire_tbl3_taylor_prod_w_vector1_range10168w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9248w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10184w(0) <= wire_tbl3_taylor_prod_w_vector1_range10179w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10178w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10185w(0) <= wire_tbl3_taylor_prod_w_vector1_range10179w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9258w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10195w(0) <= wire_tbl3_taylor_prod_w_vector1_range10190w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10189w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10196w(0) <= wire_tbl3_taylor_prod_w_vector1_range10190w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9268w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10206w(0) <= wire_tbl3_taylor_prod_w_vector1_range10201w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10200w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10207w(0) <= wire_tbl3_taylor_prod_w_vector1_range10201w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9278w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10008w(0) <= wire_tbl3_taylor_prod_w_vector1_range10003w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10002w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10009w(0) <= wire_tbl3_taylor_prod_w_vector1_range10003w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9098w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10217w(0) <= wire_tbl3_taylor_prod_w_vector1_range10212w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10211w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10218w(0) <= wire_tbl3_taylor_prod_w_vector1_range10212w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9288w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10228w(0) <= wire_tbl3_taylor_prod_w_vector1_range10223w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10222w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10229w(0) <= wire_tbl3_taylor_prod_w_vector1_range10223w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9298w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10239w(0) <= wire_tbl3_taylor_prod_w_vector1_range10234w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10233w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10240w(0) <= wire_tbl3_taylor_prod_w_vector1_range10234w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9308w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10250w(0) <= wire_tbl3_taylor_prod_w_vector1_range10245w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10244w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10251w(0) <= wire_tbl3_taylor_prod_w_vector1_range10245w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9318w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10261w(0) <= wire_tbl3_taylor_prod_w_vector1_range10256w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10255w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10262w(0) <= wire_tbl3_taylor_prod_w_vector1_range10256w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9328w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10272w(0) <= wire_tbl3_taylor_prod_w_vector1_range10267w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10266w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10273w(0) <= wire_tbl3_taylor_prod_w_vector1_range10267w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9338w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10283w(0) <= wire_tbl3_taylor_prod_w_vector1_range10278w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10277w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10284w(0) <= wire_tbl3_taylor_prod_w_vector1_range10278w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9348w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10294w(0) <= wire_tbl3_taylor_prod_w_vector1_range10289w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10288w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10295w(0) <= wire_tbl3_taylor_prod_w_vector1_range10289w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9358w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10305w(0) <= wire_tbl3_taylor_prod_w_vector1_range10300w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10299w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10306w(0) <= wire_tbl3_taylor_prod_w_vector1_range10300w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9368w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10316w(0) <= wire_tbl3_taylor_prod_w_vector1_range10311w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10310w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10317w(0) <= wire_tbl3_taylor_prod_w_vector1_range10311w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9378w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10019w(0) <= wire_tbl3_taylor_prod_w_vector1_range10014w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10013w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10020w(0) <= wire_tbl3_taylor_prod_w_vector1_range10014w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9108w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10327w(0) <= wire_tbl3_taylor_prod_w_vector1_range10322w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10321w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10328w(0) <= wire_tbl3_taylor_prod_w_vector1_range10322w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9388w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10338w(0) <= wire_tbl3_taylor_prod_w_vector1_range10333w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10332w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10339w(0) <= wire_tbl3_taylor_prod_w_vector1_range10333w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9398w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10349w(0) <= wire_tbl3_taylor_prod_w_vector1_range10344w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10343w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10350w(0) <= wire_tbl3_taylor_prod_w_vector1_range10344w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9408w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10360w(0) <= wire_tbl3_taylor_prod_w_vector1_range10355w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10354w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10361w(0) <= wire_tbl3_taylor_prod_w_vector1_range10355w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9418w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10371w(0) <= wire_tbl3_taylor_prod_w_vector1_range10366w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10365w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10372w(0) <= wire_tbl3_taylor_prod_w_vector1_range10366w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9428w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10382w(0) <= wire_tbl3_taylor_prod_w_vector1_range10377w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10376w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10383w(0) <= wire_tbl3_taylor_prod_w_vector1_range10377w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9438w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10393w(0) <= wire_tbl3_taylor_prod_w_vector1_range10388w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10387w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10394w(0) <= wire_tbl3_taylor_prod_w_vector1_range10388w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9448w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10404w(0) <= wire_tbl3_taylor_prod_w_vector1_range10399w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10398w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10405w(0) <= wire_tbl3_taylor_prod_w_vector1_range10399w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9458w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10415w(0) <= wire_tbl3_taylor_prod_w_vector1_range10410w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10409w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10416w(0) <= wire_tbl3_taylor_prod_w_vector1_range10410w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9468w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10426w(0) <= wire_tbl3_taylor_prod_w_vector1_range10421w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10420w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10427w(0) <= wire_tbl3_taylor_prod_w_vector1_range10421w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9478w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10030w(0) <= wire_tbl3_taylor_prod_w_vector1_range10025w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10024w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10031w(0) <= wire_tbl3_taylor_prod_w_vector1_range10025w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9118w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10437w(0) <= wire_tbl3_taylor_prod_w_vector1_range10432w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10431w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10438w(0) <= wire_tbl3_taylor_prod_w_vector1_range10432w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9488w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10448w(0) <= wire_tbl3_taylor_prod_w_vector1_range10443w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10442w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10449w(0) <= wire_tbl3_taylor_prod_w_vector1_range10443w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9498w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10459w(0) <= wire_tbl3_taylor_prod_w_vector1_range10454w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10453w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10460w(0) <= wire_tbl3_taylor_prod_w_vector1_range10454w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9508w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10470w(0) <= wire_tbl3_taylor_prod_w_vector1_range10465w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10464w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10471w(0) <= wire_tbl3_taylor_prod_w_vector1_range10465w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9518w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10481w(0) <= wire_tbl3_taylor_prod_w_vector1_range10476w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10475w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10482w(0) <= wire_tbl3_taylor_prod_w_vector1_range10476w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9528w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10492w(0) <= wire_tbl3_taylor_prod_w_vector1_range10487w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10486w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10493w(0) <= wire_tbl3_taylor_prod_w_vector1_range10487w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9538w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10503w(0) <= wire_tbl3_taylor_prod_w_vector1_range10498w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10497w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10504w(0) <= wire_tbl3_taylor_prod_w_vector1_range10498w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9548w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10514w(0) <= wire_tbl3_taylor_prod_w_vector1_range10509w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10508w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10515w(0) <= wire_tbl3_taylor_prod_w_vector1_range10509w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9558w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10525w(0) <= wire_tbl3_taylor_prod_w_vector1_range10520w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10519w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10526w(0) <= wire_tbl3_taylor_prod_w_vector1_range10520w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9568w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10536w(0) <= wire_tbl3_taylor_prod_w_vector1_range10531w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10530w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10537w(0) <= wire_tbl3_taylor_prod_w_vector1_range10531w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9578w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10041w(0) <= wire_tbl3_taylor_prod_w_vector1_range10036w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10035w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10042w(0) <= wire_tbl3_taylor_prod_w_vector1_range10036w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9128w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10547w(0) <= wire_tbl3_taylor_prod_w_vector1_range10542w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10541w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10548w(0) <= wire_tbl3_taylor_prod_w_vector1_range10542w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9588w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10558w(0) <= wire_tbl3_taylor_prod_w_vector1_range10553w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10552w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10559w(0) <= wire_tbl3_taylor_prod_w_vector1_range10553w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9598w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10569w(0) <= wire_tbl3_taylor_prod_w_vector1_range10564w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10563w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10570w(0) <= wire_tbl3_taylor_prod_w_vector1_range10564w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9608w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10580w(0) <= wire_tbl3_taylor_prod_w_vector1_range10575w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10574w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10581w(0) <= wire_tbl3_taylor_prod_w_vector1_range10575w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9618w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10591w(0) <= wire_tbl3_taylor_prod_w_vector1_range10586w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10585w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10592w(0) <= wire_tbl3_taylor_prod_w_vector1_range10586w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9628w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10602w(0) <= wire_tbl3_taylor_prod_w_vector1_range10597w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10596w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10603w(0) <= wire_tbl3_taylor_prod_w_vector1_range10597w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9638w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10613w(0) <= wire_tbl3_taylor_prod_w_vector1_range10608w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10607w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10614w(0) <= wire_tbl3_taylor_prod_w_vector1_range10608w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9648w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10624w(0) <= wire_tbl3_taylor_prod_w_vector1_range10619w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10618w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10625w(0) <= wire_tbl3_taylor_prod_w_vector1_range10619w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9658w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10635w(0) <= wire_tbl3_taylor_prod_w_vector1_range10630w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10629w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10636w(0) <= wire_tbl3_taylor_prod_w_vector1_range10630w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9668w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10646w(0) <= wire_tbl3_taylor_prod_w_vector1_range10641w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10640w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10647w(0) <= wire_tbl3_taylor_prod_w_vector1_range10641w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9678w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10052w(0) <= wire_tbl3_taylor_prod_w_vector1_range10047w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10046w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10053w(0) <= wire_tbl3_taylor_prod_w_vector1_range10047w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9138w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10657w(0) <= wire_tbl3_taylor_prod_w_vector1_range10652w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10651w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10658w(0) <= wire_tbl3_taylor_prod_w_vector1_range10652w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9688w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10668w(0) <= wire_tbl3_taylor_prod_w_vector1_range10663w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10662w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10669w(0) <= wire_tbl3_taylor_prod_w_vector1_range10663w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9698w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10679w(0) <= wire_tbl3_taylor_prod_w_vector1_range10674w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10673w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10680w(0) <= wire_tbl3_taylor_prod_w_vector1_range10674w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9708w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10690w(0) <= wire_tbl3_taylor_prod_w_vector1_range10685w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10684w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10691w(0) <= wire_tbl3_taylor_prod_w_vector1_range10685w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9718w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10701w(0) <= wire_tbl3_taylor_prod_w_vector1_range10696w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10695w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10702w(0) <= wire_tbl3_taylor_prod_w_vector1_range10696w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9728w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10712w(0) <= wire_tbl3_taylor_prod_w_vector1_range10707w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10706w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10713w(0) <= wire_tbl3_taylor_prod_w_vector1_range10707w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9738w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10723w(0) <= wire_tbl3_taylor_prod_w_vector1_range10718w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10717w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10724w(0) <= wire_tbl3_taylor_prod_w_vector1_range10718w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9748w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10734w(0) <= wire_tbl3_taylor_prod_w_vector1_range10729w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10728w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10735w(0) <= wire_tbl3_taylor_prod_w_vector1_range10729w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9758w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10745w(0) <= wire_tbl3_taylor_prod_w_vector1_range10740w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10739w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10746w(0) <= wire_tbl3_taylor_prod_w_vector1_range10740w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9768w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10756w(0) <= wire_tbl3_taylor_prod_w_vector1_range10751w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10750w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10757w(0) <= wire_tbl3_taylor_prod_w_vector1_range10751w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9778w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10063w(0) <= wire_tbl3_taylor_prod_w_vector1_range10058w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10057w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10064w(0) <= wire_tbl3_taylor_prod_w_vector1_range10058w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9148w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10767w(0) <= wire_tbl3_taylor_prod_w_vector1_range10762w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10761w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10768w(0) <= wire_tbl3_taylor_prod_w_vector1_range10762w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9788w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10778w(0) <= wire_tbl3_taylor_prod_w_vector1_range10773w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10772w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10779w(0) <= wire_tbl3_taylor_prod_w_vector1_range10773w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9798w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10789w(0) <= wire_tbl3_taylor_prod_w_vector1_range10784w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10783w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10790w(0) <= wire_tbl3_taylor_prod_w_vector1_range10784w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9808w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10800w(0) <= wire_tbl3_taylor_prod_w_vector1_range10795w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10794w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10801w(0) <= wire_tbl3_taylor_prod_w_vector1_range10795w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9818w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10811w(0) <= wire_tbl3_taylor_prod_w_vector1_range10806w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10805w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10812w(0) <= wire_tbl3_taylor_prod_w_vector1_range10806w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9828w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10822w(0) <= wire_tbl3_taylor_prod_w_vector1_range10817w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10816w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10823w(0) <= wire_tbl3_taylor_prod_w_vector1_range10817w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9838w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10833w(0) <= wire_tbl3_taylor_prod_w_vector1_range10828w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10827w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10834w(0) <= wire_tbl3_taylor_prod_w_vector1_range10828w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9848w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10844w(0) <= wire_tbl3_taylor_prod_w_vector1_range10839w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10838w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10845w(0) <= wire_tbl3_taylor_prod_w_vector1_range10839w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9858w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10855w(0) <= wire_tbl3_taylor_prod_w_vector1_range10850w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10849w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10856w(0) <= wire_tbl3_taylor_prod_w_vector1_range10850w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9868w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10866w(0) <= wire_tbl3_taylor_prod_w_vector1_range10861w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10860w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10867w(0) <= wire_tbl3_taylor_prod_w_vector1_range10861w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9878w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10074w(0) <= wire_tbl3_taylor_prod_w_vector1_range10069w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10068w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10075w(0) <= wire_tbl3_taylor_prod_w_vector1_range10069w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9158w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10877w(0) <= wire_tbl3_taylor_prod_w_vector1_range10872w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10871w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10878w(0) <= wire_tbl3_taylor_prod_w_vector1_range10872w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9888w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10888w(0) <= wire_tbl3_taylor_prod_w_vector1_range10883w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10882w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10889w(0) <= wire_tbl3_taylor_prod_w_vector1_range10883w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9898w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10899w(0) <= wire_tbl3_taylor_prod_w_vector1_range10894w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10893w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10900w(0) <= wire_tbl3_taylor_prod_w_vector1_range10894w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9908w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10910w(0) <= wire_tbl3_taylor_prod_w_vector1_range10905w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10904w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10911w(0) <= wire_tbl3_taylor_prod_w_vector1_range10905w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9918w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10921w(0) <= wire_tbl3_taylor_prod_w_vector1_range10916w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10915w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10922w(0) <= wire_tbl3_taylor_prod_w_vector1_range10916w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9928w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10932w(0) <= wire_tbl3_taylor_prod_w_vector1_range10927w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10926w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10933w(0) <= wire_tbl3_taylor_prod_w_vector1_range10927w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9938w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10943w(0) <= wire_tbl3_taylor_prod_w_vector1_range10938w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10937w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10944w(0) <= wire_tbl3_taylor_prod_w_vector1_range10938w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9948w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10954w(0) <= wire_tbl3_taylor_prod_w_vector1_range10949w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10948w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10955w(0) <= wire_tbl3_taylor_prod_w_vector1_range10949w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9958w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10965w(0) <= wire_tbl3_taylor_prod_w_vector1_range10960w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10959w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10966w(0) <= wire_tbl3_taylor_prod_w_vector1_range10960w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9968w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10976w(0) <= wire_tbl3_taylor_prod_w_vector1_range10971w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10970w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10977w(0) <= wire_tbl3_taylor_prod_w_vector1_range10971w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9978w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10085w(0) <= wire_tbl3_taylor_prod_w_vector1_range10080w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10079w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10086w(0) <= wire_tbl3_taylor_prod_w_vector1_range10080w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9168w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10096w(0) <= wire_tbl3_taylor_prod_w_vector1_range10091w(0) AND wire_tbl3_taylor_prod_w_car_one_adj_range10090w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10097w(0) <= wire_tbl3_taylor_prod_w_vector1_range10091w(0) AND wire_tbl3_taylor_prod_w_sum_one_range9178w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9089w(0) <= wire_tbl3_taylor_prod_w_vector2_range9083w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9082w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9090w(0) <= wire_tbl3_taylor_prod_w_vector2_range9083w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9079w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9190w(0) <= wire_tbl3_taylor_prod_w_vector2_range9185w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9022w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9191w(0) <= wire_tbl3_taylor_prod_w_vector2_range9185w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9019w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9200w(0) <= wire_tbl3_taylor_prod_w_vector2_range9195w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9016w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9201w(0) <= wire_tbl3_taylor_prod_w_vector2_range9195w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9013w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9210w(0) <= wire_tbl3_taylor_prod_w_vector2_range9205w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9010w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9211w(0) <= wire_tbl3_taylor_prod_w_vector2_range9205w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9007w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9220w(0) <= wire_tbl3_taylor_prod_w_vector2_range9215w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9004w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9221w(0) <= wire_tbl3_taylor_prod_w_vector2_range9215w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9001w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9230w(0) <= wire_tbl3_taylor_prod_w_vector2_range9225w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8998w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9231w(0) <= wire_tbl3_taylor_prod_w_vector2_range9225w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8995w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9240w(0) <= wire_tbl3_taylor_prod_w_vector2_range9235w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8992w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9241w(0) <= wire_tbl3_taylor_prod_w_vector2_range9235w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8989w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9250w(0) <= wire_tbl3_taylor_prod_w_vector2_range9245w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8986w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9251w(0) <= wire_tbl3_taylor_prod_w_vector2_range9245w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8983w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9260w(0) <= wire_tbl3_taylor_prod_w_vector2_range9255w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8980w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9261w(0) <= wire_tbl3_taylor_prod_w_vector2_range9255w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8977w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9270w(0) <= wire_tbl3_taylor_prod_w_vector2_range9265w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8974w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9271w(0) <= wire_tbl3_taylor_prod_w_vector2_range9265w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8971w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9280w(0) <= wire_tbl3_taylor_prod_w_vector2_range9275w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8968w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9281w(0) <= wire_tbl3_taylor_prod_w_vector2_range9275w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8965w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9100w(0) <= wire_tbl3_taylor_prod_w_vector2_range9095w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9076w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9101w(0) <= wire_tbl3_taylor_prod_w_vector2_range9095w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9073w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9290w(0) <= wire_tbl3_taylor_prod_w_vector2_range9285w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8962w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9291w(0) <= wire_tbl3_taylor_prod_w_vector2_range9285w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8959w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9300w(0) <= wire_tbl3_taylor_prod_w_vector2_range9295w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8956w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9301w(0) <= wire_tbl3_taylor_prod_w_vector2_range9295w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8953w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9310w(0) <= wire_tbl3_taylor_prod_w_vector2_range9305w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8950w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9311w(0) <= wire_tbl3_taylor_prod_w_vector2_range9305w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8947w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9320w(0) <= wire_tbl3_taylor_prod_w_vector2_range9315w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8944w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9321w(0) <= wire_tbl3_taylor_prod_w_vector2_range9315w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8941w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9330w(0) <= wire_tbl3_taylor_prod_w_vector2_range9325w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8938w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9331w(0) <= wire_tbl3_taylor_prod_w_vector2_range9325w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8935w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9340w(0) <= wire_tbl3_taylor_prod_w_vector2_range9335w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8932w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9341w(0) <= wire_tbl3_taylor_prod_w_vector2_range9335w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8929w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9350w(0) <= wire_tbl3_taylor_prod_w_vector2_range9345w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8926w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9351w(0) <= wire_tbl3_taylor_prod_w_vector2_range9345w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8923w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9360w(0) <= wire_tbl3_taylor_prod_w_vector2_range9355w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8920w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9361w(0) <= wire_tbl3_taylor_prod_w_vector2_range9355w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8917w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9370w(0) <= wire_tbl3_taylor_prod_w_vector2_range9365w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8914w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9371w(0) <= wire_tbl3_taylor_prod_w_vector2_range9365w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8911w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9380w(0) <= wire_tbl3_taylor_prod_w_vector2_range9375w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8908w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9381w(0) <= wire_tbl3_taylor_prod_w_vector2_range9375w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8905w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9110w(0) <= wire_tbl3_taylor_prod_w_vector2_range9105w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9070w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9111w(0) <= wire_tbl3_taylor_prod_w_vector2_range9105w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9067w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9390w(0) <= wire_tbl3_taylor_prod_w_vector2_range9385w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8902w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9391w(0) <= wire_tbl3_taylor_prod_w_vector2_range9385w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8899w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9400w(0) <= wire_tbl3_taylor_prod_w_vector2_range9395w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8896w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9401w(0) <= wire_tbl3_taylor_prod_w_vector2_range9395w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8893w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9410w(0) <= wire_tbl3_taylor_prod_w_vector2_range9405w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8890w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9411w(0) <= wire_tbl3_taylor_prod_w_vector2_range9405w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8887w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9420w(0) <= wire_tbl3_taylor_prod_w_vector2_range9415w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8884w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9421w(0) <= wire_tbl3_taylor_prod_w_vector2_range9415w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8881w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9430w(0) <= wire_tbl3_taylor_prod_w_vector2_range9425w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8878w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9431w(0) <= wire_tbl3_taylor_prod_w_vector2_range9425w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8875w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9440w(0) <= wire_tbl3_taylor_prod_w_vector2_range9435w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8872w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9441w(0) <= wire_tbl3_taylor_prod_w_vector2_range9435w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8869w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9450w(0) <= wire_tbl3_taylor_prod_w_vector2_range9445w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8866w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9451w(0) <= wire_tbl3_taylor_prod_w_vector2_range9445w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8863w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9460w(0) <= wire_tbl3_taylor_prod_w_vector2_range9455w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8860w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9461w(0) <= wire_tbl3_taylor_prod_w_vector2_range9455w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8857w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9470w(0) <= wire_tbl3_taylor_prod_w_vector2_range9465w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8854w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9471w(0) <= wire_tbl3_taylor_prod_w_vector2_range9465w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8851w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9480w(0) <= wire_tbl3_taylor_prod_w_vector2_range9475w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8848w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9481w(0) <= wire_tbl3_taylor_prod_w_vector2_range9475w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8845w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9120w(0) <= wire_tbl3_taylor_prod_w_vector2_range9115w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9064w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9121w(0) <= wire_tbl3_taylor_prod_w_vector2_range9115w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9061w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9490w(0) <= wire_tbl3_taylor_prod_w_vector2_range9485w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8842w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9491w(0) <= wire_tbl3_taylor_prod_w_vector2_range9485w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8839w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9500w(0) <= wire_tbl3_taylor_prod_w_vector2_range9495w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8836w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9501w(0) <= wire_tbl3_taylor_prod_w_vector2_range9495w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8833w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9510w(0) <= wire_tbl3_taylor_prod_w_vector2_range9505w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8830w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9511w(0) <= wire_tbl3_taylor_prod_w_vector2_range9505w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8827w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9520w(0) <= wire_tbl3_taylor_prod_w_vector2_range9515w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8824w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9521w(0) <= wire_tbl3_taylor_prod_w_vector2_range9515w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8821w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9530w(0) <= wire_tbl3_taylor_prod_w_vector2_range9525w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8818w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9531w(0) <= wire_tbl3_taylor_prod_w_vector2_range9525w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8815w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9540w(0) <= wire_tbl3_taylor_prod_w_vector2_range9535w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8812w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9541w(0) <= wire_tbl3_taylor_prod_w_vector2_range9535w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8809w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9550w(0) <= wire_tbl3_taylor_prod_w_vector2_range9545w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8806w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9551w(0) <= wire_tbl3_taylor_prod_w_vector2_range9545w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8803w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9560w(0) <= wire_tbl3_taylor_prod_w_vector2_range9555w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8800w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9561w(0) <= wire_tbl3_taylor_prod_w_vector2_range9555w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8797w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9570w(0) <= wire_tbl3_taylor_prod_w_vector2_range9565w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8794w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9571w(0) <= wire_tbl3_taylor_prod_w_vector2_range9565w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8791w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9580w(0) <= wire_tbl3_taylor_prod_w_vector2_range9575w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8788w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9581w(0) <= wire_tbl3_taylor_prod_w_vector2_range9575w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8785w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9130w(0) <= wire_tbl3_taylor_prod_w_vector2_range9125w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9058w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9131w(0) <= wire_tbl3_taylor_prod_w_vector2_range9125w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9055w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9590w(0) <= wire_tbl3_taylor_prod_w_vector2_range9585w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8782w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9591w(0) <= wire_tbl3_taylor_prod_w_vector2_range9585w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8779w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9600w(0) <= wire_tbl3_taylor_prod_w_vector2_range9595w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8776w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9601w(0) <= wire_tbl3_taylor_prod_w_vector2_range9595w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8773w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9610w(0) <= wire_tbl3_taylor_prod_w_vector2_range9605w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8770w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9611w(0) <= wire_tbl3_taylor_prod_w_vector2_range9605w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8767w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9620w(0) <= wire_tbl3_taylor_prod_w_vector2_range9615w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8764w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9621w(0) <= wire_tbl3_taylor_prod_w_vector2_range9615w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8761w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9630w(0) <= wire_tbl3_taylor_prod_w_vector2_range9625w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8758w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9631w(0) <= wire_tbl3_taylor_prod_w_vector2_range9625w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8755w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9640w(0) <= wire_tbl3_taylor_prod_w_vector2_range9635w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8752w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9641w(0) <= wire_tbl3_taylor_prod_w_vector2_range9635w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8749w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9650w(0) <= wire_tbl3_taylor_prod_w_vector2_range9645w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8746w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9651w(0) <= wire_tbl3_taylor_prod_w_vector2_range9645w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8743w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9660w(0) <= wire_tbl3_taylor_prod_w_vector2_range9655w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8740w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9661w(0) <= wire_tbl3_taylor_prod_w_vector2_range9655w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8737w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9670w(0) <= wire_tbl3_taylor_prod_w_vector2_range9665w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8734w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9671w(0) <= wire_tbl3_taylor_prod_w_vector2_range9665w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8731w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9680w(0) <= wire_tbl3_taylor_prod_w_vector2_range9675w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8728w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9681w(0) <= wire_tbl3_taylor_prod_w_vector2_range9675w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8724w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9140w(0) <= wire_tbl3_taylor_prod_w_vector2_range9135w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9052w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9141w(0) <= wire_tbl3_taylor_prod_w_vector2_range9135w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9049w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9690w(0) <= wire_tbl3_taylor_prod_w_vector2_range9685w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8723w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9691w(0) <= wire_tbl3_taylor_prod_w_vector2_range9685w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8719w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9700w(0) <= wire_tbl3_taylor_prod_w_vector2_range9695w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8718w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9701w(0) <= wire_tbl3_taylor_prod_w_vector2_range9695w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8714w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9710w(0) <= wire_tbl3_taylor_prod_w_vector2_range9705w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8712w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9711w(0) <= wire_tbl3_taylor_prod_w_vector2_range9705w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8710w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9720w(0) <= wire_tbl3_taylor_prod_w_vector2_range9715w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8708w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9721w(0) <= wire_tbl3_taylor_prod_w_vector2_range9715w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8706w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9730w(0) <= wire_tbl3_taylor_prod_w_vector2_range9725w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8704w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9731w(0) <= wire_tbl3_taylor_prod_w_vector2_range9725w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8702w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9740w(0) <= wire_tbl3_taylor_prod_w_vector2_range9735w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8700w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9741w(0) <= wire_tbl3_taylor_prod_w_vector2_range9735w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8698w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9750w(0) <= wire_tbl3_taylor_prod_w_vector2_range9745w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8696w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9751w(0) <= wire_tbl3_taylor_prod_w_vector2_range9745w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8694w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9760w(0) <= wire_tbl3_taylor_prod_w_vector2_range9755w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8692w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9761w(0) <= wire_tbl3_taylor_prod_w_vector2_range9755w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8690w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9770w(0) <= wire_tbl3_taylor_prod_w_vector2_range9765w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8688w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9771w(0) <= wire_tbl3_taylor_prod_w_vector2_range9765w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8686w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9780w(0) <= wire_tbl3_taylor_prod_w_vector2_range9775w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8684w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9781w(0) <= wire_tbl3_taylor_prod_w_vector2_range9775w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8682w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9150w(0) <= wire_tbl3_taylor_prod_w_vector2_range9145w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9046w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9151w(0) <= wire_tbl3_taylor_prod_w_vector2_range9145w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9043w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9790w(0) <= wire_tbl3_taylor_prod_w_vector2_range9785w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8680w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9791w(0) <= wire_tbl3_taylor_prod_w_vector2_range9785w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8678w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9800w(0) <= wire_tbl3_taylor_prod_w_vector2_range9795w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8676w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9801w(0) <= wire_tbl3_taylor_prod_w_vector2_range9795w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8674w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9810w(0) <= wire_tbl3_taylor_prod_w_vector2_range9805w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8672w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9811w(0) <= wire_tbl3_taylor_prod_w_vector2_range9805w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8670w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9820w(0) <= wire_tbl3_taylor_prod_w_vector2_range9815w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8668w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9821w(0) <= wire_tbl3_taylor_prod_w_vector2_range9815w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8666w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9830w(0) <= wire_tbl3_taylor_prod_w_vector2_range9825w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8664w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9831w(0) <= wire_tbl3_taylor_prod_w_vector2_range9825w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8662w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9840w(0) <= wire_tbl3_taylor_prod_w_vector2_range9835w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8660w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9841w(0) <= wire_tbl3_taylor_prod_w_vector2_range9835w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8658w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9850w(0) <= wire_tbl3_taylor_prod_w_vector2_range9845w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8656w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9851w(0) <= wire_tbl3_taylor_prod_w_vector2_range9845w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8654w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9860w(0) <= wire_tbl3_taylor_prod_w_vector2_range9855w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8652w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9861w(0) <= wire_tbl3_taylor_prod_w_vector2_range9855w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8650w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9870w(0) <= wire_tbl3_taylor_prod_w_vector2_range9865w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8648w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9871w(0) <= wire_tbl3_taylor_prod_w_vector2_range9865w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8646w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9880w(0) <= wire_tbl3_taylor_prod_w_vector2_range9875w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8644w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9881w(0) <= wire_tbl3_taylor_prod_w_vector2_range9875w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8642w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9160w(0) <= wire_tbl3_taylor_prod_w_vector2_range9155w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9040w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9161w(0) <= wire_tbl3_taylor_prod_w_vector2_range9155w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9037w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9890w(0) <= wire_tbl3_taylor_prod_w_vector2_range9885w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8640w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9891w(0) <= wire_tbl3_taylor_prod_w_vector2_range9885w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8638w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9900w(0) <= wire_tbl3_taylor_prod_w_vector2_range9895w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8636w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9901w(0) <= wire_tbl3_taylor_prod_w_vector2_range9895w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8634w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9910w(0) <= wire_tbl3_taylor_prod_w_vector2_range9905w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8632w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9911w(0) <= wire_tbl3_taylor_prod_w_vector2_range9905w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8630w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9920w(0) <= wire_tbl3_taylor_prod_w_vector2_range9915w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8628w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9921w(0) <= wire_tbl3_taylor_prod_w_vector2_range9915w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8626w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9930w(0) <= wire_tbl3_taylor_prod_w_vector2_range9925w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8624w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9931w(0) <= wire_tbl3_taylor_prod_w_vector2_range9925w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8622w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9940w(0) <= wire_tbl3_taylor_prod_w_vector2_range9935w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8620w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9941w(0) <= wire_tbl3_taylor_prod_w_vector2_range9935w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8618w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9950w(0) <= wire_tbl3_taylor_prod_w_vector2_range9945w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8616w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9951w(0) <= wire_tbl3_taylor_prod_w_vector2_range9945w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8614w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9960w(0) <= wire_tbl3_taylor_prod_w_vector2_range9955w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8612w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9961w(0) <= wire_tbl3_taylor_prod_w_vector2_range9955w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8610w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9970w(0) <= wire_tbl3_taylor_prod_w_vector2_range9965w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8608w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9971w(0) <= wire_tbl3_taylor_prod_w_vector2_range9965w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8606w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9980w(0) <= wire_tbl3_taylor_prod_w_vector2_range9975w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range8603w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9981w(0) <= wire_tbl3_taylor_prod_w_vector2_range9975w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range8600w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9170w(0) <= wire_tbl3_taylor_prod_w_vector2_range9165w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9034w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9171w(0) <= wire_tbl3_taylor_prod_w_vector2_range9165w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9031w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9180w(0) <= wire_tbl3_taylor_prod_w_vector2_range9175w(0) AND wire_tbl3_taylor_prod_w_neg_lsb_range9028w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9181w(0) <= wire_tbl3_taylor_prod_w_vector2_range9175w(0) AND wire_tbl3_taylor_prod_w_neg_msb_range9025w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9080w9081w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9080w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9020w9021w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9020w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9014w9015w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9014w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9008w9009w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9008w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9002w9003w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9002w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8996w8997w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8996w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8990w8991w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8990w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8984w8985w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8984w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8978w8979w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8978w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8972w8973w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8972w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8966w8967w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8966w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9074w9075w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9074w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8960w8961w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8960w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8954w8955w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8954w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8948w8949w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8948w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8942w8943w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8942w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8936w8937w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8936w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8930w8931w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8930w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8924w8925w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8924w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8918w8919w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8918w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8912w8913w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8912w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8906w8907w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8906w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9068w9069w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9068w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8900w8901w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8900w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8894w8895w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8894w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8888w8889w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8888w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8882w8883w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8882w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8876w8877w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8876w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8870w8871w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8870w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8864w8865w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8864w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8858w8859w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8858w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8852w8853w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8852w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8846w8847w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8846w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9062w9063w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9062w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8840w8841w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8840w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8834w8835w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8834w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8828w8829w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8828w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8822w8823w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8822w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8816w8817w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8816w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8810w8811w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8810w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8804w8805w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8804w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8798w8799w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8798w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8792w8793w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8792w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8786w8787w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8786w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9056w9057w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9056w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8780w8781w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8780w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8774w8775w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8774w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8768w8769w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8768w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8762w8763w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8762w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8756w8757w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8756w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8750w8751w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8750w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8744w8745w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8744w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8738w8739w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8738w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8732w8733w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8732w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8726w8727w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8726w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9050w9051w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9050w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8721w8722w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8721w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8716w8717w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range8716w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9044w9045w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9044w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9038w9039w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9038w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9032w9033w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9032w(0);
	wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9026w9027w(0) <= NOT wire_tbl3_taylor_prod_w_lsb_prod_wo_range9026w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9077w9078w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9077w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9017w9018w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9017w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9011w9012w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9011w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9005w9006w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9005w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8999w9000w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8999w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8993w8994w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8993w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8987w8988w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8987w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8981w8982w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8981w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8975w8976w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8975w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8969w8970w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8969w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8963w8964w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8963w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9071w9072w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9071w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8957w8958w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8957w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8951w8952w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8951w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8945w8946w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8945w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8939w8940w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8939w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8933w8934w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8933w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8927w8928w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8927w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8921w8922w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8921w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8915w8916w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8915w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8909w8910w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8909w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8903w8904w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8903w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9065w9066w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9065w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8897w8898w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8897w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8891w8892w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8891w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8885w8886w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8885w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8879w8880w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8879w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8873w8874w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8873w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8867w8868w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8867w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8861w8862w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8861w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8855w8856w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8855w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8849w8850w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8849w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8843w8844w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8843w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9059w9060w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9059w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8837w8838w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8837w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8831w8832w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8831w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8825w8826w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8825w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8819w8820w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8819w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8813w8814w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8813w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8807w8808w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8807w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8801w8802w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8801w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8795w8796w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8795w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8789w8790w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8789w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8783w8784w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8783w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9053w9054w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9053w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8777w8778w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8777w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8771w8772w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8771w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8765w8766w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8765w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8759w8760w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8759w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8753w8754w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8753w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8747w8748w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8747w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8741w8742w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8741w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8735w8736w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8735w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8729w8730w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range8729w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9047w9048w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9047w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9041w9042w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9041w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9035w9036w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9035w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9029w9030w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9029w(0);
	wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9023w9024w(0) <= NOT wire_tbl3_taylor_prod_w_msb_prod_wo_range9023w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range9990w9997w9998w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9997w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9996w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10102w10108w10109w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10108w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10107w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10113w10119w10120w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10119w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10118w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10124w10130w10131w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10130w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10129w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10135w10141w10142w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10141w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10140w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10146w10152w10153w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10152w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10151w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10157w10163w10164w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10163w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10162w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10168w10174w10175w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10174w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10173w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10179w10185w10186w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10185w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10184w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10190w10196w10197w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10196w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10195w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10201w10207w10208w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10207w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10206w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10003w10009w10010w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10009w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10008w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10212w10218w10219w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10218w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10217w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10223w10229w10230w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10229w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10228w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10234w10240w10241w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10240w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10239w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10245w10251w10252w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10251w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10250w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10256w10262w10263w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10262w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10261w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10267w10273w10274w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10273w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10272w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10278w10284w10285w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10284w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10283w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10289w10295w10296w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10295w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10294w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10300w10306w10307w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10306w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10305w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10311w10317w10318w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10317w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10316w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10014w10020w10021w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10020w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10019w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10322w10328w10329w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10328w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10327w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10333w10339w10340w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10339w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10338w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10344w10350w10351w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10350w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10349w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10355w10361w10362w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10361w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10360w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10366w10372w10373w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10372w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10371w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10377w10383w10384w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10383w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10382w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10388w10394w10395w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10394w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10393w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10399w10405w10406w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10405w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10404w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10410w10416w10417w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10416w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10415w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10421w10427w10428w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10427w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10426w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10025w10031w10032w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10031w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10030w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10432w10438w10439w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10438w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10437w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10443w10449w10450w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10449w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10448w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10454w10460w10461w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10460w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10459w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10465w10471w10472w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10471w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10470w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10476w10482w10483w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10482w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10481w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10487w10493w10494w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10493w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10492w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10498w10504w10505w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10504w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10503w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10509w10515w10516w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10515w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10514w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10520w10526w10527w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10526w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10525w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10531w10537w10538w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10537w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10536w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10036w10042w10043w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10042w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10041w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10542w10548w10549w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10548w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10547w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10553w10559w10560w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10559w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10558w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10564w10570w10571w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10570w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10569w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10575w10581w10582w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10581w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10580w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10586w10592w10593w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10592w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10591w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10597w10603w10604w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10603w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10602w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10608w10614w10615w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10614w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10613w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10619w10625w10626w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10625w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10624w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10630w10636w10637w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10636w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10635w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10641w10647w10648w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10647w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10646w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10047w10053w10054w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10053w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10052w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10652w10658w10659w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10658w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10657w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10663w10669w10670w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10669w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10668w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10674w10680w10681w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10680w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10679w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10685w10691w10692w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10691w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10690w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10696w10702w10703w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10702w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10701w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10707w10713w10714w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10713w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10712w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10718w10724w10725w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10724w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10723w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10729w10735w10736w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10735w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10734w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10740w10746w10747w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10746w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10745w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10751w10757w10758w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10757w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10756w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10058w10064w10065w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10064w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10063w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10762w10768w10769w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10768w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10767w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10773w10779w10780w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10779w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10778w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10784w10790w10791w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10790w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10789w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10795w10801w10802w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10801w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10800w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10806w10812w10813w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10812w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10811w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10817w10823w10824w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10823w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10822w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10828w10834w10835w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10834w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10833w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10839w10845w10846w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10845w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10844w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10850w10856w10857w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10856w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10855w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10861w10867w10868w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10867w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10866w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10069w10075w10076w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10075w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10074w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10872w10878w10879w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10878w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10877w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10883w10889w10890w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10889w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10888w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10894w10900w10901w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10900w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10899w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10905w10911w10912w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10911w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10910w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10916w10922w10923w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10922w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10921w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10927w10933w10934w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10933w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10932w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10938w10944w10945w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10944w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10943w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10949w10955w10956w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10955w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10954w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10960w10966w10967w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10966w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10965w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10971w10977w10978w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10977w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10976w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10080w10086w10087w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10086w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10085w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10091w10097w10098w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10097w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10096w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9083w9090w9091w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9090w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9089w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9185w9191w9192w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9191w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9190w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9195w9201w9202w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9201w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9200w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9205w9211w9212w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9211w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9210w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9215w9221w9222w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9221w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9220w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9225w9231w9232w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9231w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9230w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9235w9241w9242w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9241w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9240w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9245w9251w9252w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9251w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9250w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9255w9261w9262w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9261w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9260w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9265w9271w9272w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9271w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9270w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9275w9281w9282w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9281w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9280w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9095w9101w9102w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9101w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9100w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9285w9291w9292w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9291w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9290w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9295w9301w9302w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9301w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9300w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9305w9311w9312w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9311w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9310w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9315w9321w9322w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9321w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9320w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9325w9331w9332w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9331w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9330w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9335w9341w9342w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9341w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9340w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9345w9351w9352w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9351w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9350w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9355w9361w9362w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9361w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9360w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9365w9371w9372w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9371w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9370w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9375w9381w9382w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9381w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9380w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9105w9111w9112w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9111w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9110w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9385w9391w9392w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9391w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9390w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9395w9401w9402w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9401w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9400w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9405w9411w9412w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9411w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9410w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9415w9421w9422w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9421w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9420w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9425w9431w9432w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9431w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9430w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9435w9441w9442w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9441w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9440w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9445w9451w9452w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9451w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9450w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9455w9461w9462w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9461w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9460w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9465w9471w9472w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9471w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9470w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9475w9481w9482w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9481w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9480w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9115w9121w9122w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9121w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9120w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9485w9491w9492w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9491w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9490w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9495w9501w9502w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9501w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9500w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9505w9511w9512w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9511w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9510w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9515w9521w9522w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9521w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9520w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9525w9531w9532w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9531w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9530w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9535w9541w9542w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9541w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9540w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9545w9551w9552w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9551w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9550w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9555w9561w9562w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9561w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9560w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9565w9571w9572w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9571w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9570w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9575w9581w9582w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9581w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9580w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9125w9131w9132w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9131w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9130w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9585w9591w9592w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9591w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9590w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9595w9601w9602w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9601w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9600w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9605w9611w9612w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9611w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9610w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9615w9621w9622w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9621w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9620w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9625w9631w9632w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9631w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9630w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9635w9641w9642w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9641w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9640w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9645w9651w9652w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9651w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9650w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9655w9661w9662w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9661w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9660w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9665w9671w9672w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9671w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9670w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9675w9681w9682w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9681w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9680w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9135w9141w9142w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9141w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9140w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9685w9691w9692w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9691w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9690w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9695w9701w9702w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9701w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9700w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9705w9711w9712w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9711w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9710w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9715w9721w9722w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9721w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9720w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9725w9731w9732w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9731w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9730w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9735w9741w9742w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9741w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9740w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9745w9751w9752w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9751w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9750w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9755w9761w9762w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9761w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9760w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9765w9771w9772w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9771w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9770w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9775w9781w9782w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9781w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9780w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9145w9151w9152w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9151w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9150w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9785w9791w9792w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9791w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9790w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9795w9801w9802w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9801w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9800w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9805w9811w9812w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9811w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9810w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9815w9821w9822w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9821w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9820w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9825w9831w9832w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9831w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9830w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9835w9841w9842w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9841w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9840w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9845w9851w9852w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9851w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9850w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9855w9861w9862w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9861w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9860w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9865w9871w9872w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9871w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9870w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9875w9881w9882w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9881w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9880w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9155w9161w9162w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9161w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9160w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9885w9891w9892w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9891w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9890w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9895w9901w9902w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9901w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9900w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9905w9911w9912w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9911w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9910w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9915w9921w9922w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9921w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9920w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9925w9931w9932w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9931w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9930w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9935w9941w9942w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9941w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9940w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9945w9951w9952w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9951w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9950w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9955w9961w9962w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9961w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9960w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9965w9971w9972w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9971w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9970w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9975w9981w9982w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9981w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9980w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9165w9171w9172w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9171w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9170w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9175w9181w9182w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9181w(0) OR wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9180w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector1_range9990w9997w9998w9999w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range9990w9997w9998w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9086w9995w(0);
	wire_tbl3_taylor_prod_w10110w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10102w10108w10109w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9188w10106w(0);
	wire_tbl3_taylor_prod_w10121w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10113w10119w10120w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9198w10117w(0);
	wire_tbl3_taylor_prod_w10132w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10124w10130w10131w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9208w10128w(0);
	wire_tbl3_taylor_prod_w10143w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10135w10141w10142w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9218w10139w(0);
	wire_tbl3_taylor_prod_w10154w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10146w10152w10153w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9228w10150w(0);
	wire_tbl3_taylor_prod_w10165w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10157w10163w10164w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9238w10161w(0);
	wire_tbl3_taylor_prod_w10176w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10168w10174w10175w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9248w10172w(0);
	wire_tbl3_taylor_prod_w10187w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10179w10185w10186w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9258w10183w(0);
	wire_tbl3_taylor_prod_w10198w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10190w10196w10197w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9268w10194w(0);
	wire_tbl3_taylor_prod_w10209w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10201w10207w10208w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9278w10205w(0);
	wire_tbl3_taylor_prod_w10011w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10003w10009w10010w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9098w10007w(0);
	wire_tbl3_taylor_prod_w10220w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10212w10218w10219w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9288w10216w(0);
	wire_tbl3_taylor_prod_w10231w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10223w10229w10230w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9298w10227w(0);
	wire_tbl3_taylor_prod_w10242w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10234w10240w10241w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9308w10238w(0);
	wire_tbl3_taylor_prod_w10253w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10245w10251w10252w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9318w10249w(0);
	wire_tbl3_taylor_prod_w10264w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10256w10262w10263w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9328w10260w(0);
	wire_tbl3_taylor_prod_w10275w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10267w10273w10274w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9338w10271w(0);
	wire_tbl3_taylor_prod_w10286w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10278w10284w10285w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9348w10282w(0);
	wire_tbl3_taylor_prod_w10297w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10289w10295w10296w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9358w10293w(0);
	wire_tbl3_taylor_prod_w10308w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10300w10306w10307w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9368w10304w(0);
	wire_tbl3_taylor_prod_w10319w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10311w10317w10318w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9378w10315w(0);
	wire_tbl3_taylor_prod_w10022w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10014w10020w10021w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9108w10018w(0);
	wire_tbl3_taylor_prod_w10330w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10322w10328w10329w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9388w10326w(0);
	wire_tbl3_taylor_prod_w10341w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10333w10339w10340w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9398w10337w(0);
	wire_tbl3_taylor_prod_w10352w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10344w10350w10351w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9408w10348w(0);
	wire_tbl3_taylor_prod_w10363w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10355w10361w10362w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9418w10359w(0);
	wire_tbl3_taylor_prod_w10374w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10366w10372w10373w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9428w10370w(0);
	wire_tbl3_taylor_prod_w10385w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10377w10383w10384w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9438w10381w(0);
	wire_tbl3_taylor_prod_w10396w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10388w10394w10395w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9448w10392w(0);
	wire_tbl3_taylor_prod_w10407w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10399w10405w10406w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9458w10403w(0);
	wire_tbl3_taylor_prod_w10418w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10410w10416w10417w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9468w10414w(0);
	wire_tbl3_taylor_prod_w10429w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10421w10427w10428w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9478w10425w(0);
	wire_tbl3_taylor_prod_w10033w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10025w10031w10032w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9118w10029w(0);
	wire_tbl3_taylor_prod_w10440w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10432w10438w10439w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9488w10436w(0);
	wire_tbl3_taylor_prod_w10451w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10443w10449w10450w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9498w10447w(0);
	wire_tbl3_taylor_prod_w10462w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10454w10460w10461w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9508w10458w(0);
	wire_tbl3_taylor_prod_w10473w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10465w10471w10472w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9518w10469w(0);
	wire_tbl3_taylor_prod_w10484w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10476w10482w10483w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9528w10480w(0);
	wire_tbl3_taylor_prod_w10495w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10487w10493w10494w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9538w10491w(0);
	wire_tbl3_taylor_prod_w10506w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10498w10504w10505w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9548w10502w(0);
	wire_tbl3_taylor_prod_w10517w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10509w10515w10516w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9558w10513w(0);
	wire_tbl3_taylor_prod_w10528w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10520w10526w10527w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9568w10524w(0);
	wire_tbl3_taylor_prod_w10539w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10531w10537w10538w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9578w10535w(0);
	wire_tbl3_taylor_prod_w10044w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10036w10042w10043w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9128w10040w(0);
	wire_tbl3_taylor_prod_w10550w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10542w10548w10549w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9588w10546w(0);
	wire_tbl3_taylor_prod_w10561w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10553w10559w10560w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9598w10557w(0);
	wire_tbl3_taylor_prod_w10572w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10564w10570w10571w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9608w10568w(0);
	wire_tbl3_taylor_prod_w10583w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10575w10581w10582w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9618w10579w(0);
	wire_tbl3_taylor_prod_w10594w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10586w10592w10593w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9628w10590w(0);
	wire_tbl3_taylor_prod_w10605w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10597w10603w10604w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9638w10601w(0);
	wire_tbl3_taylor_prod_w10616w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10608w10614w10615w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9648w10612w(0);
	wire_tbl3_taylor_prod_w10627w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10619w10625w10626w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9658w10623w(0);
	wire_tbl3_taylor_prod_w10638w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10630w10636w10637w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9668w10634w(0);
	wire_tbl3_taylor_prod_w10649w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10641w10647w10648w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9678w10645w(0);
	wire_tbl3_taylor_prod_w10055w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10047w10053w10054w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9138w10051w(0);
	wire_tbl3_taylor_prod_w10660w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10652w10658w10659w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9688w10656w(0);
	wire_tbl3_taylor_prod_w10671w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10663w10669w10670w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9698w10667w(0);
	wire_tbl3_taylor_prod_w10682w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10674w10680w10681w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9708w10678w(0);
	wire_tbl3_taylor_prod_w10693w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10685w10691w10692w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9718w10689w(0);
	wire_tbl3_taylor_prod_w10704w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10696w10702w10703w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9728w10700w(0);
	wire_tbl3_taylor_prod_w10715w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10707w10713w10714w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9738w10711w(0);
	wire_tbl3_taylor_prod_w10726w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10718w10724w10725w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9748w10722w(0);
	wire_tbl3_taylor_prod_w10737w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10729w10735w10736w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9758w10733w(0);
	wire_tbl3_taylor_prod_w10748w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10740w10746w10747w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9768w10744w(0);
	wire_tbl3_taylor_prod_w10759w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10751w10757w10758w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9778w10755w(0);
	wire_tbl3_taylor_prod_w10066w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10058w10064w10065w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9148w10062w(0);
	wire_tbl3_taylor_prod_w10770w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10762w10768w10769w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9788w10766w(0);
	wire_tbl3_taylor_prod_w10781w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10773w10779w10780w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9798w10777w(0);
	wire_tbl3_taylor_prod_w10792w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10784w10790w10791w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9808w10788w(0);
	wire_tbl3_taylor_prod_w10803w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10795w10801w10802w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9818w10799w(0);
	wire_tbl3_taylor_prod_w10814w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10806w10812w10813w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9828w10810w(0);
	wire_tbl3_taylor_prod_w10825w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10817w10823w10824w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9838w10821w(0);
	wire_tbl3_taylor_prod_w10836w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10828w10834w10835w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9848w10832w(0);
	wire_tbl3_taylor_prod_w10847w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10839w10845w10846w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9858w10843w(0);
	wire_tbl3_taylor_prod_w10858w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10850w10856w10857w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9868w10854w(0);
	wire_tbl3_taylor_prod_w10869w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10861w10867w10868w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9878w10865w(0);
	wire_tbl3_taylor_prod_w10077w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10069w10075w10076w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9158w10073w(0);
	wire_tbl3_taylor_prod_w10880w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10872w10878w10879w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9888w10876w(0);
	wire_tbl3_taylor_prod_w10891w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10883w10889w10890w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9898w10887w(0);
	wire_tbl3_taylor_prod_w10902w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10894w10900w10901w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9908w10898w(0);
	wire_tbl3_taylor_prod_w10913w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10905w10911w10912w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9918w10909w(0);
	wire_tbl3_taylor_prod_w10924w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10916w10922w10923w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9928w10920w(0);
	wire_tbl3_taylor_prod_w10935w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10927w10933w10934w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9938w10931w(0);
	wire_tbl3_taylor_prod_w10946w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10938w10944w10945w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9948w10942w(0);
	wire_tbl3_taylor_prod_w10957w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10949w10955w10956w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9958w10953w(0);
	wire_tbl3_taylor_prod_w10968w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10960w10966w10967w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9968w10964w(0);
	wire_tbl3_taylor_prod_w10979w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10971w10977w10978w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9978w10975w(0);
	wire_tbl3_taylor_prod_w10088w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10080w10086w10087w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9168w10084w(0);
	wire_tbl3_taylor_prod_w10099w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10091w10097w10098w(0) OR wire_tbl3_taylor_prod_w_lg_w_sum_one_range9178w10095w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9083w9090w9091w9092w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9083w9090w9091w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9079w9088w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9185w9191w9192w9193w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9185w9191w9192w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9019w9189w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9195w9201w9202w9203w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9195w9201w9202w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9013w9199w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9205w9211w9212w9213w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9205w9211w9212w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9007w9209w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9215w9221w9222w9223w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9215w9221w9222w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9001w9219w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9225w9231w9232w9233w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9225w9231w9232w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8995w9229w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9235w9241w9242w9243w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9235w9241w9242w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8989w9239w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9245w9251w9252w9253w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9245w9251w9252w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8983w9249w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9255w9261w9262w9263w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9255w9261w9262w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8977w9259w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9265w9271w9272w9273w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9265w9271w9272w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8971w9269w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9275w9281w9282w9283w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9275w9281w9282w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8965w9279w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9095w9101w9102w9103w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9095w9101w9102w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9073w9099w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9285w9291w9292w9293w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9285w9291w9292w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8959w9289w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9295w9301w9302w9303w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9295w9301w9302w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8953w9299w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9305w9311w9312w9313w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9305w9311w9312w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8947w9309w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9315w9321w9322w9323w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9315w9321w9322w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8941w9319w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9325w9331w9332w9333w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9325w9331w9332w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8935w9329w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9335w9341w9342w9343w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9335w9341w9342w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8929w9339w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9345w9351w9352w9353w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9345w9351w9352w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8923w9349w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9355w9361w9362w9363w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9355w9361w9362w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8917w9359w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9365w9371w9372w9373w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9365w9371w9372w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8911w9369w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9375w9381w9382w9383w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9375w9381w9382w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8905w9379w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9105w9111w9112w9113w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9105w9111w9112w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9067w9109w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9385w9391w9392w9393w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9385w9391w9392w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8899w9389w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9395w9401w9402w9403w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9395w9401w9402w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8893w9399w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9405w9411w9412w9413w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9405w9411w9412w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8887w9409w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9415w9421w9422w9423w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9415w9421w9422w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8881w9419w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9425w9431w9432w9433w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9425w9431w9432w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8875w9429w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9435w9441w9442w9443w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9435w9441w9442w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8869w9439w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9445w9451w9452w9453w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9445w9451w9452w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8863w9449w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9455w9461w9462w9463w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9455w9461w9462w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8857w9459w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9465w9471w9472w9473w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9465w9471w9472w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8851w9469w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9475w9481w9482w9483w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9475w9481w9482w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8845w9479w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9115w9121w9122w9123w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9115w9121w9122w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9061w9119w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9485w9491w9492w9493w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9485w9491w9492w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8839w9489w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9495w9501w9502w9503w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9495w9501w9502w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8833w9499w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9505w9511w9512w9513w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9505w9511w9512w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8827w9509w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9515w9521w9522w9523w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9515w9521w9522w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8821w9519w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9525w9531w9532w9533w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9525w9531w9532w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8815w9529w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9535w9541w9542w9543w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9535w9541w9542w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8809w9539w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9545w9551w9552w9553w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9545w9551w9552w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8803w9549w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9555w9561w9562w9563w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9555w9561w9562w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8797w9559w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9565w9571w9572w9573w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9565w9571w9572w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8791w9569w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9575w9581w9582w9583w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9575w9581w9582w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8785w9579w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9125w9131w9132w9133w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9125w9131w9132w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9055w9129w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9585w9591w9592w9593w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9585w9591w9592w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8779w9589w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9595w9601w9602w9603w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9595w9601w9602w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8773w9599w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9605w9611w9612w9613w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9605w9611w9612w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8767w9609w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9615w9621w9622w9623w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9615w9621w9622w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8761w9619w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9625w9631w9632w9633w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9625w9631w9632w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8755w9629w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9635w9641w9642w9643w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9635w9641w9642w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8749w9639w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9645w9651w9652w9653w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9645w9651w9652w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8743w9649w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9655w9661w9662w9663w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9655w9661w9662w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8737w9659w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9665w9671w9672w9673w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9665w9671w9672w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8731w9669w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9675w9681w9682w9683w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9675w9681w9682w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8724w9679w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9135w9141w9142w9143w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9135w9141w9142w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9049w9139w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9685w9691w9692w9693w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9685w9691w9692w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8719w9689w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9695w9701w9702w9703w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9695w9701w9702w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8714w9699w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9705w9711w9712w9713w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9705w9711w9712w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8710w9709w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9715w9721w9722w9723w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9715w9721w9722w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8706w9719w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9725w9731w9732w9733w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9725w9731w9732w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8702w9729w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9735w9741w9742w9743w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9735w9741w9742w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8698w9739w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9745w9751w9752w9753w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9745w9751w9752w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8694w9749w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9755w9761w9762w9763w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9755w9761w9762w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8690w9759w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9765w9771w9772w9773w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9765w9771w9772w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8686w9769w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9775w9781w9782w9783w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9775w9781w9782w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8682w9779w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9145w9151w9152w9153w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9145w9151w9152w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9043w9149w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9785w9791w9792w9793w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9785w9791w9792w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8678w9789w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9795w9801w9802w9803w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9795w9801w9802w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8674w9799w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9805w9811w9812w9813w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9805w9811w9812w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8670w9809w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9815w9821w9822w9823w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9815w9821w9822w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8666w9819w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9825w9831w9832w9833w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9825w9831w9832w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8662w9829w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9835w9841w9842w9843w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9835w9841w9842w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8658w9839w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9845w9851w9852w9853w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9845w9851w9852w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8654w9849w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9855w9861w9862w9863w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9855w9861w9862w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8650w9859w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9865w9871w9872w9873w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9865w9871w9872w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8646w9869w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9875w9881w9882w9883w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9875w9881w9882w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8642w9879w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9155w9161w9162w9163w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9155w9161w9162w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9037w9159w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9885w9891w9892w9893w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9885w9891w9892w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8638w9889w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9895w9901w9902w9903w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9895w9901w9902w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8634w9899w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9905w9911w9912w9913w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9905w9911w9912w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8630w9909w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9915w9921w9922w9923w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9915w9921w9922w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8626w9919w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9925w9931w9932w9933w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9925w9931w9932w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8622w9929w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9935w9941w9942w9943w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9935w9941w9942w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8618w9939w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9945w9951w9952w9953w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9945w9951w9952w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8614w9949w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9955w9961w9962w9963w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9955w9961w9962w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8610w9959w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9965w9971w9972w9973w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9965w9971w9972w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8606w9969w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9975w9981w9982w9983w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9975w9981w9982w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range8600w9979w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9165w9171w9172w9173w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9165w9171w9172w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9031w9169w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9175w9181w9182w9183w(0) <= wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9175w9181w9182w(0) OR wire_tbl3_taylor_prod_w_lg_w_neg_msb_range9025w9179w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range9990w9991w9992w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9991w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range9988w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10102w10103w10104w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10103w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10101w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10113w10114w10115w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10114w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10112w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10124w10125w10126w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10125w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10123w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10135w10136w10137w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10136w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10134w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10146w10147w10148w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10147w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10145w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10157w10158w10159w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10158w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10156w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10168w10169w10170w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10169w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10167w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10179w10180w10181w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10180w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10178w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10190w10191w10192w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10191w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10189w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10201w10202w10203w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10202w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10200w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10003w10004w10005w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10004w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10002w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10212w10213w10214w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10213w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10211w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10223w10224w10225w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10224w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10222w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10234w10235w10236w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10235w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10233w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10245w10246w10247w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10246w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10244w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10256w10257w10258w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10257w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10255w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10267w10268w10269w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10268w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10266w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10278w10279w10280w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10279w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10277w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10289w10290w10291w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10290w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10288w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10300w10301w10302w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10301w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10299w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10311w10312w10313w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10312w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10310w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10014w10015w10016w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10015w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10013w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10322w10323w10324w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10323w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10321w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10333w10334w10335w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10334w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10332w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10344w10345w10346w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10345w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10343w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10355w10356w10357w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10356w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10354w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10366w10367w10368w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10367w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10365w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10377w10378w10379w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10378w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10376w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10388w10389w10390w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10389w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10387w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10399w10400w10401w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10400w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10398w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10410w10411w10412w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10411w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10409w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10421w10422w10423w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10422w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10420w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10025w10026w10027w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10026w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10024w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10432w10433w10434w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10433w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10431w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10443w10444w10445w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10444w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10442w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10454w10455w10456w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10455w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10453w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10465w10466w10467w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10466w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10464w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10476w10477w10478w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10477w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10475w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10487w10488w10489w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10488w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10486w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10498w10499w10500w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10499w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10497w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10509w10510w10511w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10510w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10508w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10520w10521w10522w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10521w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10519w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10531w10532w10533w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10532w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10530w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10036w10037w10038w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10037w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10035w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10542w10543w10544w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10543w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10541w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10553w10554w10555w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10554w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10552w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10564w10565w10566w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10565w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10563w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10575w10576w10577w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10576w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10574w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10586w10587w10588w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10587w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10585w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10597w10598w10599w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10598w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10596w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10608w10609w10610w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10609w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10607w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10619w10620w10621w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10620w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10618w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10630w10631w10632w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10631w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10629w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10641w10642w10643w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10642w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10640w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10047w10048w10049w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10048w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10046w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10652w10653w10654w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10653w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10651w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10663w10664w10665w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10664w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10662w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10674w10675w10676w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10675w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10673w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10685w10686w10687w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10686w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10684w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10696w10697w10698w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10697w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10695w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10707w10708w10709w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10708w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10706w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10718w10719w10720w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10719w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10717w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10729w10730w10731w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10730w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10728w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10740w10741w10742w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10741w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10739w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10751w10752w10753w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10752w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10750w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10058w10059w10060w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10059w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10057w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10762w10763w10764w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10763w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10761w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10773w10774w10775w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10774w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10772w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10784w10785w10786w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10785w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10783w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10795w10796w10797w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10796w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10794w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10806w10807w10808w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10807w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10805w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10817w10818w10819w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10818w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10816w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10828w10829w10830w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10829w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10827w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10839w10840w10841w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10840w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10838w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10850w10851w10852w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10851w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10849w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10861w10862w10863w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10862w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10860w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10069w10070w10071w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10070w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10068w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10872w10873w10874w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10873w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10871w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10883w10884w10885w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10884w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10882w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10894w10895w10896w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10895w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10893w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10905w10906w10907w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10906w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10904w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10916w10917w10918w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10917w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10915w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10927w10928w10929w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10928w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10926w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10938w10939w10940w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10939w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10937w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10949w10950w10951w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10950w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10948w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10960w10961w10962w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10961w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10959w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10971w10972w10973w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10972w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10970w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10080w10081w10082w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10081w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10079w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10091w10092w10093w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10092w(0) XOR wire_tbl3_taylor_prod_w_car_one_adj_range10090w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9083w9084w9085w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9084w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9082w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9185w9186w9187w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9186w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9022w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9195w9196w9197w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9196w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9016w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9205w9206w9207w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9206w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9010w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9215w9216w9217w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9216w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9004w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9225w9226w9227w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9226w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8998w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9235w9236w9237w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9236w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8992w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9245w9246w9247w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9246w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8986w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9255w9256w9257w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9256w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8980w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9265w9266w9267w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9266w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8974w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9275w9276w9277w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9276w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8968w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9095w9096w9097w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9096w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9076w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9285w9286w9287w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9286w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8962w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9295w9296w9297w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9296w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8956w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9305w9306w9307w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9306w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8950w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9315w9316w9317w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9316w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8944w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9325w9326w9327w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9326w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8938w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9335w9336w9337w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9336w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8932w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9345w9346w9347w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9346w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8926w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9355w9356w9357w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9356w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8920w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9365w9366w9367w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9366w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8914w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9375w9376w9377w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9376w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8908w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9105w9106w9107w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9106w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9070w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9385w9386w9387w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9386w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8902w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9395w9396w9397w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9396w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8896w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9405w9406w9407w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9406w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8890w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9415w9416w9417w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9416w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8884w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9425w9426w9427w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9426w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8878w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9435w9436w9437w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9436w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8872w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9445w9446w9447w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9446w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8866w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9455w9456w9457w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9456w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8860w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9465w9466w9467w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9466w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8854w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9475w9476w9477w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9476w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8848w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9115w9116w9117w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9116w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9064w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9485w9486w9487w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9486w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8842w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9495w9496w9497w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9496w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8836w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9505w9506w9507w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9506w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8830w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9515w9516w9517w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9516w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8824w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9525w9526w9527w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9526w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8818w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9535w9536w9537w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9536w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8812w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9545w9546w9547w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9546w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8806w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9555w9556w9557w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9556w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8800w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9565w9566w9567w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9566w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8794w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9575w9576w9577w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9576w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8788w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9125w9126w9127w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9126w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9058w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9585w9586w9587w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9586w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8782w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9595w9596w9597w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9596w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8776w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9605w9606w9607w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9606w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8770w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9615w9616w9617w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9616w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8764w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9625w9626w9627w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9626w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8758w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9635w9636w9637w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9636w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8752w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9645w9646w9647w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9646w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8746w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9655w9656w9657w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9656w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8740w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9665w9666w9667w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9666w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8734w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9675w9676w9677w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9676w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8728w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9135w9136w9137w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9136w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9052w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9685w9686w9687w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9686w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8723w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9695w9696w9697w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9696w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8718w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9705w9706w9707w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9706w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8712w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9715w9716w9717w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9716w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8708w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9725w9726w9727w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9726w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8704w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9735w9736w9737w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9736w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8700w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9745w9746w9747w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9746w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8696w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9755w9756w9757w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9756w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8692w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9765w9766w9767w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9766w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8688w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9775w9776w9777w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9776w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8684w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9145w9146w9147w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9146w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9046w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9785w9786w9787w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9786w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8680w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9795w9796w9797w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9796w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8676w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9805w9806w9807w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9806w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8672w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9815w9816w9817w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9816w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8668w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9825w9826w9827w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9826w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8664w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9835w9836w9837w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9836w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8660w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9845w9846w9847w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9846w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8656w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9855w9856w9857w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9856w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8652w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9865w9866w9867w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9866w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8648w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9875w9876w9877w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9876w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8644w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9155w9156w9157w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9156w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9040w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9885w9886w9887w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9886w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8640w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9895w9896w9897w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9896w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8636w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9905w9906w9907w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9906w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8632w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9915w9916w9917w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9916w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8628w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9925w9926w9927w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9926w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8624w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9935w9936w9937w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9936w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8620w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9945w9946w9947w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9946w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8616w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9955w9956w9957w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9956w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8612w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9965w9966w9967w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9966w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8608w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9975w9976w9977w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9976w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range8603w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9165w9166w9167w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9166w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9034w(0);
	wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9175w9176w9177w(0) <= wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9176w(0) XOR wire_tbl3_taylor_prod_w_neg_lsb_range9028w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range9990w9991w(0) <= wire_tbl3_taylor_prod_w_vector1_range9990w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9086w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10102w10103w(0) <= wire_tbl3_taylor_prod_w_vector1_range10102w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9188w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10113w10114w(0) <= wire_tbl3_taylor_prod_w_vector1_range10113w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9198w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10124w10125w(0) <= wire_tbl3_taylor_prod_w_vector1_range10124w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9208w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10135w10136w(0) <= wire_tbl3_taylor_prod_w_vector1_range10135w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9218w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10146w10147w(0) <= wire_tbl3_taylor_prod_w_vector1_range10146w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9228w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10157w10158w(0) <= wire_tbl3_taylor_prod_w_vector1_range10157w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9238w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10168w10169w(0) <= wire_tbl3_taylor_prod_w_vector1_range10168w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9248w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10179w10180w(0) <= wire_tbl3_taylor_prod_w_vector1_range10179w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9258w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10190w10191w(0) <= wire_tbl3_taylor_prod_w_vector1_range10190w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9268w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10201w10202w(0) <= wire_tbl3_taylor_prod_w_vector1_range10201w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9278w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10003w10004w(0) <= wire_tbl3_taylor_prod_w_vector1_range10003w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9098w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10212w10213w(0) <= wire_tbl3_taylor_prod_w_vector1_range10212w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9288w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10223w10224w(0) <= wire_tbl3_taylor_prod_w_vector1_range10223w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9298w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10234w10235w(0) <= wire_tbl3_taylor_prod_w_vector1_range10234w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9308w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10245w10246w(0) <= wire_tbl3_taylor_prod_w_vector1_range10245w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9318w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10256w10257w(0) <= wire_tbl3_taylor_prod_w_vector1_range10256w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9328w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10267w10268w(0) <= wire_tbl3_taylor_prod_w_vector1_range10267w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9338w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10278w10279w(0) <= wire_tbl3_taylor_prod_w_vector1_range10278w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9348w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10289w10290w(0) <= wire_tbl3_taylor_prod_w_vector1_range10289w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9358w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10300w10301w(0) <= wire_tbl3_taylor_prod_w_vector1_range10300w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9368w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10311w10312w(0) <= wire_tbl3_taylor_prod_w_vector1_range10311w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9378w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10014w10015w(0) <= wire_tbl3_taylor_prod_w_vector1_range10014w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9108w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10322w10323w(0) <= wire_tbl3_taylor_prod_w_vector1_range10322w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9388w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10333w10334w(0) <= wire_tbl3_taylor_prod_w_vector1_range10333w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9398w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10344w10345w(0) <= wire_tbl3_taylor_prod_w_vector1_range10344w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9408w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10355w10356w(0) <= wire_tbl3_taylor_prod_w_vector1_range10355w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9418w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10366w10367w(0) <= wire_tbl3_taylor_prod_w_vector1_range10366w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9428w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10377w10378w(0) <= wire_tbl3_taylor_prod_w_vector1_range10377w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9438w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10388w10389w(0) <= wire_tbl3_taylor_prod_w_vector1_range10388w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9448w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10399w10400w(0) <= wire_tbl3_taylor_prod_w_vector1_range10399w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9458w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10410w10411w(0) <= wire_tbl3_taylor_prod_w_vector1_range10410w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9468w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10421w10422w(0) <= wire_tbl3_taylor_prod_w_vector1_range10421w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9478w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10025w10026w(0) <= wire_tbl3_taylor_prod_w_vector1_range10025w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9118w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10432w10433w(0) <= wire_tbl3_taylor_prod_w_vector1_range10432w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9488w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10443w10444w(0) <= wire_tbl3_taylor_prod_w_vector1_range10443w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9498w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10454w10455w(0) <= wire_tbl3_taylor_prod_w_vector1_range10454w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9508w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10465w10466w(0) <= wire_tbl3_taylor_prod_w_vector1_range10465w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9518w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10476w10477w(0) <= wire_tbl3_taylor_prod_w_vector1_range10476w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9528w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10487w10488w(0) <= wire_tbl3_taylor_prod_w_vector1_range10487w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9538w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10498w10499w(0) <= wire_tbl3_taylor_prod_w_vector1_range10498w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9548w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10509w10510w(0) <= wire_tbl3_taylor_prod_w_vector1_range10509w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9558w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10520w10521w(0) <= wire_tbl3_taylor_prod_w_vector1_range10520w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9568w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10531w10532w(0) <= wire_tbl3_taylor_prod_w_vector1_range10531w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9578w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10036w10037w(0) <= wire_tbl3_taylor_prod_w_vector1_range10036w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9128w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10542w10543w(0) <= wire_tbl3_taylor_prod_w_vector1_range10542w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9588w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10553w10554w(0) <= wire_tbl3_taylor_prod_w_vector1_range10553w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9598w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10564w10565w(0) <= wire_tbl3_taylor_prod_w_vector1_range10564w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9608w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10575w10576w(0) <= wire_tbl3_taylor_prod_w_vector1_range10575w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9618w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10586w10587w(0) <= wire_tbl3_taylor_prod_w_vector1_range10586w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9628w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10597w10598w(0) <= wire_tbl3_taylor_prod_w_vector1_range10597w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9638w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10608w10609w(0) <= wire_tbl3_taylor_prod_w_vector1_range10608w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9648w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10619w10620w(0) <= wire_tbl3_taylor_prod_w_vector1_range10619w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9658w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10630w10631w(0) <= wire_tbl3_taylor_prod_w_vector1_range10630w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9668w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10641w10642w(0) <= wire_tbl3_taylor_prod_w_vector1_range10641w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9678w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10047w10048w(0) <= wire_tbl3_taylor_prod_w_vector1_range10047w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9138w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10652w10653w(0) <= wire_tbl3_taylor_prod_w_vector1_range10652w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9688w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10663w10664w(0) <= wire_tbl3_taylor_prod_w_vector1_range10663w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9698w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10674w10675w(0) <= wire_tbl3_taylor_prod_w_vector1_range10674w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9708w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10685w10686w(0) <= wire_tbl3_taylor_prod_w_vector1_range10685w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9718w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10696w10697w(0) <= wire_tbl3_taylor_prod_w_vector1_range10696w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9728w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10707w10708w(0) <= wire_tbl3_taylor_prod_w_vector1_range10707w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9738w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10718w10719w(0) <= wire_tbl3_taylor_prod_w_vector1_range10718w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9748w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10729w10730w(0) <= wire_tbl3_taylor_prod_w_vector1_range10729w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9758w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10740w10741w(0) <= wire_tbl3_taylor_prod_w_vector1_range10740w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9768w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10751w10752w(0) <= wire_tbl3_taylor_prod_w_vector1_range10751w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9778w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10058w10059w(0) <= wire_tbl3_taylor_prod_w_vector1_range10058w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9148w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10762w10763w(0) <= wire_tbl3_taylor_prod_w_vector1_range10762w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9788w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10773w10774w(0) <= wire_tbl3_taylor_prod_w_vector1_range10773w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9798w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10784w10785w(0) <= wire_tbl3_taylor_prod_w_vector1_range10784w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9808w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10795w10796w(0) <= wire_tbl3_taylor_prod_w_vector1_range10795w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9818w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10806w10807w(0) <= wire_tbl3_taylor_prod_w_vector1_range10806w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9828w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10817w10818w(0) <= wire_tbl3_taylor_prod_w_vector1_range10817w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9838w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10828w10829w(0) <= wire_tbl3_taylor_prod_w_vector1_range10828w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9848w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10839w10840w(0) <= wire_tbl3_taylor_prod_w_vector1_range10839w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9858w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10850w10851w(0) <= wire_tbl3_taylor_prod_w_vector1_range10850w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9868w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10861w10862w(0) <= wire_tbl3_taylor_prod_w_vector1_range10861w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9878w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10069w10070w(0) <= wire_tbl3_taylor_prod_w_vector1_range10069w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9158w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10872w10873w(0) <= wire_tbl3_taylor_prod_w_vector1_range10872w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9888w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10883w10884w(0) <= wire_tbl3_taylor_prod_w_vector1_range10883w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9898w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10894w10895w(0) <= wire_tbl3_taylor_prod_w_vector1_range10894w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9908w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10905w10906w(0) <= wire_tbl3_taylor_prod_w_vector1_range10905w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9918w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10916w10917w(0) <= wire_tbl3_taylor_prod_w_vector1_range10916w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9928w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10927w10928w(0) <= wire_tbl3_taylor_prod_w_vector1_range10927w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9938w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10938w10939w(0) <= wire_tbl3_taylor_prod_w_vector1_range10938w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9948w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10949w10950w(0) <= wire_tbl3_taylor_prod_w_vector1_range10949w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9958w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10960w10961w(0) <= wire_tbl3_taylor_prod_w_vector1_range10960w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9968w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10971w10972w(0) <= wire_tbl3_taylor_prod_w_vector1_range10971w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9978w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10080w10081w(0) <= wire_tbl3_taylor_prod_w_vector1_range10080w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9168w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector1_range10091w10092w(0) <= wire_tbl3_taylor_prod_w_vector1_range10091w(0) XOR wire_tbl3_taylor_prod_w_sum_one_range9178w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9083w9084w(0) <= wire_tbl3_taylor_prod_w_vector2_range9083w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9079w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9185w9186w(0) <= wire_tbl3_taylor_prod_w_vector2_range9185w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9019w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9195w9196w(0) <= wire_tbl3_taylor_prod_w_vector2_range9195w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9013w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9205w9206w(0) <= wire_tbl3_taylor_prod_w_vector2_range9205w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9007w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9215w9216w(0) <= wire_tbl3_taylor_prod_w_vector2_range9215w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9001w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9225w9226w(0) <= wire_tbl3_taylor_prod_w_vector2_range9225w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8995w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9235w9236w(0) <= wire_tbl3_taylor_prod_w_vector2_range9235w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8989w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9245w9246w(0) <= wire_tbl3_taylor_prod_w_vector2_range9245w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8983w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9255w9256w(0) <= wire_tbl3_taylor_prod_w_vector2_range9255w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8977w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9265w9266w(0) <= wire_tbl3_taylor_prod_w_vector2_range9265w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8971w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9275w9276w(0) <= wire_tbl3_taylor_prod_w_vector2_range9275w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8965w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9095w9096w(0) <= wire_tbl3_taylor_prod_w_vector2_range9095w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9073w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9285w9286w(0) <= wire_tbl3_taylor_prod_w_vector2_range9285w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8959w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9295w9296w(0) <= wire_tbl3_taylor_prod_w_vector2_range9295w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8953w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9305w9306w(0) <= wire_tbl3_taylor_prod_w_vector2_range9305w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8947w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9315w9316w(0) <= wire_tbl3_taylor_prod_w_vector2_range9315w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8941w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9325w9326w(0) <= wire_tbl3_taylor_prod_w_vector2_range9325w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8935w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9335w9336w(0) <= wire_tbl3_taylor_prod_w_vector2_range9335w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8929w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9345w9346w(0) <= wire_tbl3_taylor_prod_w_vector2_range9345w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8923w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9355w9356w(0) <= wire_tbl3_taylor_prod_w_vector2_range9355w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8917w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9365w9366w(0) <= wire_tbl3_taylor_prod_w_vector2_range9365w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8911w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9375w9376w(0) <= wire_tbl3_taylor_prod_w_vector2_range9375w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8905w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9105w9106w(0) <= wire_tbl3_taylor_prod_w_vector2_range9105w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9067w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9385w9386w(0) <= wire_tbl3_taylor_prod_w_vector2_range9385w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8899w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9395w9396w(0) <= wire_tbl3_taylor_prod_w_vector2_range9395w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8893w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9405w9406w(0) <= wire_tbl3_taylor_prod_w_vector2_range9405w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8887w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9415w9416w(0) <= wire_tbl3_taylor_prod_w_vector2_range9415w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8881w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9425w9426w(0) <= wire_tbl3_taylor_prod_w_vector2_range9425w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8875w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9435w9436w(0) <= wire_tbl3_taylor_prod_w_vector2_range9435w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8869w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9445w9446w(0) <= wire_tbl3_taylor_prod_w_vector2_range9445w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8863w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9455w9456w(0) <= wire_tbl3_taylor_prod_w_vector2_range9455w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8857w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9465w9466w(0) <= wire_tbl3_taylor_prod_w_vector2_range9465w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8851w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9475w9476w(0) <= wire_tbl3_taylor_prod_w_vector2_range9475w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8845w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9115w9116w(0) <= wire_tbl3_taylor_prod_w_vector2_range9115w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9061w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9485w9486w(0) <= wire_tbl3_taylor_prod_w_vector2_range9485w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8839w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9495w9496w(0) <= wire_tbl3_taylor_prod_w_vector2_range9495w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8833w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9505w9506w(0) <= wire_tbl3_taylor_prod_w_vector2_range9505w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8827w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9515w9516w(0) <= wire_tbl3_taylor_prod_w_vector2_range9515w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8821w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9525w9526w(0) <= wire_tbl3_taylor_prod_w_vector2_range9525w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8815w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9535w9536w(0) <= wire_tbl3_taylor_prod_w_vector2_range9535w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8809w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9545w9546w(0) <= wire_tbl3_taylor_prod_w_vector2_range9545w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8803w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9555w9556w(0) <= wire_tbl3_taylor_prod_w_vector2_range9555w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8797w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9565w9566w(0) <= wire_tbl3_taylor_prod_w_vector2_range9565w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8791w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9575w9576w(0) <= wire_tbl3_taylor_prod_w_vector2_range9575w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8785w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9125w9126w(0) <= wire_tbl3_taylor_prod_w_vector2_range9125w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9055w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9585w9586w(0) <= wire_tbl3_taylor_prod_w_vector2_range9585w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8779w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9595w9596w(0) <= wire_tbl3_taylor_prod_w_vector2_range9595w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8773w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9605w9606w(0) <= wire_tbl3_taylor_prod_w_vector2_range9605w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8767w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9615w9616w(0) <= wire_tbl3_taylor_prod_w_vector2_range9615w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8761w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9625w9626w(0) <= wire_tbl3_taylor_prod_w_vector2_range9625w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8755w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9635w9636w(0) <= wire_tbl3_taylor_prod_w_vector2_range9635w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8749w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9645w9646w(0) <= wire_tbl3_taylor_prod_w_vector2_range9645w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8743w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9655w9656w(0) <= wire_tbl3_taylor_prod_w_vector2_range9655w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8737w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9665w9666w(0) <= wire_tbl3_taylor_prod_w_vector2_range9665w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8731w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9675w9676w(0) <= wire_tbl3_taylor_prod_w_vector2_range9675w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8724w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9135w9136w(0) <= wire_tbl3_taylor_prod_w_vector2_range9135w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9049w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9685w9686w(0) <= wire_tbl3_taylor_prod_w_vector2_range9685w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8719w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9695w9696w(0) <= wire_tbl3_taylor_prod_w_vector2_range9695w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8714w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9705w9706w(0) <= wire_tbl3_taylor_prod_w_vector2_range9705w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8710w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9715w9716w(0) <= wire_tbl3_taylor_prod_w_vector2_range9715w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8706w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9725w9726w(0) <= wire_tbl3_taylor_prod_w_vector2_range9725w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8702w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9735w9736w(0) <= wire_tbl3_taylor_prod_w_vector2_range9735w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8698w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9745w9746w(0) <= wire_tbl3_taylor_prod_w_vector2_range9745w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8694w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9755w9756w(0) <= wire_tbl3_taylor_prod_w_vector2_range9755w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8690w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9765w9766w(0) <= wire_tbl3_taylor_prod_w_vector2_range9765w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8686w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9775w9776w(0) <= wire_tbl3_taylor_prod_w_vector2_range9775w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8682w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9145w9146w(0) <= wire_tbl3_taylor_prod_w_vector2_range9145w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9043w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9785w9786w(0) <= wire_tbl3_taylor_prod_w_vector2_range9785w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8678w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9795w9796w(0) <= wire_tbl3_taylor_prod_w_vector2_range9795w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8674w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9805w9806w(0) <= wire_tbl3_taylor_prod_w_vector2_range9805w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8670w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9815w9816w(0) <= wire_tbl3_taylor_prod_w_vector2_range9815w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8666w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9825w9826w(0) <= wire_tbl3_taylor_prod_w_vector2_range9825w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8662w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9835w9836w(0) <= wire_tbl3_taylor_prod_w_vector2_range9835w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8658w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9845w9846w(0) <= wire_tbl3_taylor_prod_w_vector2_range9845w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8654w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9855w9856w(0) <= wire_tbl3_taylor_prod_w_vector2_range9855w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8650w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9865w9866w(0) <= wire_tbl3_taylor_prod_w_vector2_range9865w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8646w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9875w9876w(0) <= wire_tbl3_taylor_prod_w_vector2_range9875w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8642w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9155w9156w(0) <= wire_tbl3_taylor_prod_w_vector2_range9155w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9037w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9885w9886w(0) <= wire_tbl3_taylor_prod_w_vector2_range9885w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8638w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9895w9896w(0) <= wire_tbl3_taylor_prod_w_vector2_range9895w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8634w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9905w9906w(0) <= wire_tbl3_taylor_prod_w_vector2_range9905w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8630w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9915w9916w(0) <= wire_tbl3_taylor_prod_w_vector2_range9915w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8626w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9925w9926w(0) <= wire_tbl3_taylor_prod_w_vector2_range9925w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8622w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9935w9936w(0) <= wire_tbl3_taylor_prod_w_vector2_range9935w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8618w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9945w9946w(0) <= wire_tbl3_taylor_prod_w_vector2_range9945w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8614w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9955w9956w(0) <= wire_tbl3_taylor_prod_w_vector2_range9955w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8610w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9965w9966w(0) <= wire_tbl3_taylor_prod_w_vector2_range9965w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8606w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9975w9976w(0) <= wire_tbl3_taylor_prod_w_vector2_range9975w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range8600w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9165w9166w(0) <= wire_tbl3_taylor_prod_w_vector2_range9165w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9031w(0);
	wire_tbl3_taylor_prod_w_lg_w_vector2_range9175w9176w(0) <= wire_tbl3_taylor_prod_w_vector2_range9175w(0) XOR wire_tbl3_taylor_prod_w_neg_msb_range9025w(0);
	car_one <= ( wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9975w9981w9982w9983w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9965w9971w9972w9973w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9955w9961w9962w9963w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9945w9951w9952w9953w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9935w9941w9942w9943w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9925w9931w9932w9933w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9915w9921w9922w9923w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9905w9911w9912w9913w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9895w9901w9902w9903w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9885w9891w9892w9893w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9875w9881w9882w9883w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9865w9871w9872w9873w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9855w9861w9862w9863w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9845w9851w9852w9853w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9835w9841w9842w9843w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9825w9831w9832w9833w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9815w9821w9822w9823w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9805w9811w9812w9813w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9795w9801w9802w9803w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9785w9791w9792w9793w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9775w9781w9782w9783w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9765w9771w9772w9773w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9755w9761w9762w9763w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9745w9751w9752w9753w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9735w9741w9742w9743w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9725w9731w9732w9733w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9715w9721w9722w9723w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9705w9711w9712w9713w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9695w9701w9702w9703w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9685w9691w9692w9693w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9675w9681w9682w9683w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9665w9671w9672w9673w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9655w9661w9662w9663w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9645w9651w9652w9653w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9635w9641w9642w9643w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9625w9631w9632w9633w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9615w9621w9622w9623w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9605w9611w9612w9613w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9595w9601w9602w9603w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9585w9591w9592w9593w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9575w9581w9582w9583w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9565w9571w9572w9573w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9555w9561w9562w9563w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9545w9551w9552w9553w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9535w9541w9542w9543w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9525w9531w9532w9533w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9515w9521w9522w9523w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9505w9511w9512w9513w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9495w9501w9502w9503w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9485w9491w9492w9493w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9475w9481w9482w9483w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9465w9471w9472w9473w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9455w9461w9462w9463w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9445w9451w9452w9453w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9435w9441w9442w9443w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9425w9431w9432w9433w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9415w9421w9422w9423w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9405w9411w9412w9413w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9395w9401w9402w9403w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9385w9391w9392w9393w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9375w9381w9382w9383w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9365w9371w9372w9373w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9355w9361w9362w9363w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9345w9351w9352w9353w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9335w9341w9342w9343w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9325w9331w9332w9333w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9315w9321w9322w9323w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9305w9311w9312w9313w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9295w9301w9302w9303w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9285w9291w9292w9293w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9275w9281w9282w9283w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9265w9271w9272w9273w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9255w9261w9262w9263w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9245w9251w9252w9253w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9235w9241w9242w9243w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9225w9231w9232w9233w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9215w9221w9222w9223w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9205w9211w9212w9213w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9195w9201w9202w9203w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9185w9191w9192w9193w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9175w9181w9182w9183w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9165w9171w9172w9173w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9155w9161w9162w9163w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9145w9151w9152w9153w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9135w9141w9142w9143w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9125w9131w9132w9133w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9115w9121w9122w9123w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9105w9111w9112w9113w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9095w9101w9102w9103w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector2_range9083w9090w9091w9092w);
	car_one_adj <= ( car_one(88 DOWNTO 0) & "1");
	car_two <= ( wire_tbl3_taylor_prod_w10979w & wire_tbl3_taylor_prod_w10968w & wire_tbl3_taylor_prod_w10957w & wire_tbl3_taylor_prod_w10946w & wire_tbl3_taylor_prod_w10935w & wire_tbl3_taylor_prod_w10924w & wire_tbl3_taylor_prod_w10913w & wire_tbl3_taylor_prod_w10902w & wire_tbl3_taylor_prod_w10891w & wire_tbl3_taylor_prod_w10880w & wire_tbl3_taylor_prod_w10869w & wire_tbl3_taylor_prod_w10858w & wire_tbl3_taylor_prod_w10847w & wire_tbl3_taylor_prod_w10836w & wire_tbl3_taylor_prod_w10825w & wire_tbl3_taylor_prod_w10814w & wire_tbl3_taylor_prod_w10803w & wire_tbl3_taylor_prod_w10792w & wire_tbl3_taylor_prod_w10781w & wire_tbl3_taylor_prod_w10770w & wire_tbl3_taylor_prod_w10759w & wire_tbl3_taylor_prod_w10748w & wire_tbl3_taylor_prod_w10737w & wire_tbl3_taylor_prod_w10726w & wire_tbl3_taylor_prod_w10715w & wire_tbl3_taylor_prod_w10704w & wire_tbl3_taylor_prod_w10693w & wire_tbl3_taylor_prod_w10682w & wire_tbl3_taylor_prod_w10671w & wire_tbl3_taylor_prod_w10660w & wire_tbl3_taylor_prod_w10649w & wire_tbl3_taylor_prod_w10638w & wire_tbl3_taylor_prod_w10627w & wire_tbl3_taylor_prod_w10616w & wire_tbl3_taylor_prod_w10605w & wire_tbl3_taylor_prod_w10594w & wire_tbl3_taylor_prod_w10583w & wire_tbl3_taylor_prod_w10572w & wire_tbl3_taylor_prod_w10561w & wire_tbl3_taylor_prod_w10550w & wire_tbl3_taylor_prod_w10539w & wire_tbl3_taylor_prod_w10528w & wire_tbl3_taylor_prod_w10517w & wire_tbl3_taylor_prod_w10506w & wire_tbl3_taylor_prod_w10495w & wire_tbl3_taylor_prod_w10484w & wire_tbl3_taylor_prod_w10473w & wire_tbl3_taylor_prod_w10462w & wire_tbl3_taylor_prod_w10451w & wire_tbl3_taylor_prod_w10440w & wire_tbl3_taylor_prod_w10429w & wire_tbl3_taylor_prod_w10418w & wire_tbl3_taylor_prod_w10407w & wire_tbl3_taylor_prod_w10396w & wire_tbl3_taylor_prod_w10385w & wire_tbl3_taylor_prod_w10374w & wire_tbl3_taylor_prod_w10363w & wire_tbl3_taylor_prod_w10352w & wire_tbl3_taylor_prod_w10341w & wire_tbl3_taylor_prod_w10330w & wire_tbl3_taylor_prod_w10319w & wire_tbl3_taylor_prod_w10308w & wire_tbl3_taylor_prod_w10297w & wire_tbl3_taylor_prod_w10286w
 & wire_tbl3_taylor_prod_w10275w & wire_tbl3_taylor_prod_w10264w & wire_tbl3_taylor_prod_w10253w & wire_tbl3_taylor_prod_w10242w & wire_tbl3_taylor_prod_w10231w & wire_tbl3_taylor_prod_w10220w & wire_tbl3_taylor_prod_w10209w & wire_tbl3_taylor_prod_w10198w & wire_tbl3_taylor_prod_w10187w & wire_tbl3_taylor_prod_w10176w & wire_tbl3_taylor_prod_w10165w & wire_tbl3_taylor_prod_w10154w & wire_tbl3_taylor_prod_w10143w & wire_tbl3_taylor_prod_w10132w & wire_tbl3_taylor_prod_w10121w & wire_tbl3_taylor_prod_w10110w & wire_tbl3_taylor_prod_w10099w & wire_tbl3_taylor_prod_w10088w & wire_tbl3_taylor_prod_w10077w & wire_tbl3_taylor_prod_w10066w & wire_tbl3_taylor_prod_w10055w & wire_tbl3_taylor_prod_w10044w & wire_tbl3_taylor_prod_w10033w & wire_tbl3_taylor_prod_w10022w & wire_tbl3_taylor_prod_w10011w & wire_tbl3_taylor_prod_w_lg_w_lg_w_lg_w_vector1_range9990w9997w9998w9999w);
	car_two_adj <= ( car_two(88 DOWNTO 0) & "1");
	car_two_wo <= car_two_adj_reg0;
	lowest_bits_wi <= lsb_prod_wo(30 DOWNTO 0);
	lowest_bits_wo <= lowest_bits_wi_reg2;
	lsb_prod_wi <= wire_lsb_prod_result;
	lsb_prod_wo <= lsb_prod_wi_reg0;
	mid_prod_wi <= wire_mid_prod_result;
	mid_prod_wo <= mid_prod_wi_reg0;
	msb_prod_out <= wire_msb_prod_result;
	msb_prod_wi <= msb_prod_out;
	msb_prod_wo <= msb_prod_wi_reg0;
	neg_lsb <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8716w8717w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8721w8722w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8726w8727w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8732w8733w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8738w8739w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8744w8745w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8750w8751w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8756w8757w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8762w8763w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8768w8769w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8774w8775w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8780w8781w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8786w8787w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8792w8793w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8798w8799w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8804w8805w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8810w8811w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8816w8817w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8822w8823w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8828w8829w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8834w8835w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8840w8841w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8846w8847w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8852w8853w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8858w8859w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8864w8865w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8870w8871w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8876w8877w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8882w8883w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8888w8889w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8894w8895w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8900w8901w
 & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8906w8907w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8912w8913w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8918w8919w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8924w8925w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8930w8931w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8936w8937w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8942w8943w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8948w8949w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8954w8955w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8960w8961w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8966w8967w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8972w8973w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8978w8979w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8984w8985w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8990w8991w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range8996w8997w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9002w9003w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9008w9009w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9014w9015w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9020w9021w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9026w9027w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9032w9033w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9038w9039w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9044w9045w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9050w9051w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9056w9057w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9062w9063w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9068w9069w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9074w9075w & wire_tbl3_taylor_prod_w_lg_w_lsb_prod_wo_range9080w9081w);
	neg_msb <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8729w8730w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8735w8736w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8741w8742w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8747w8748w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8753w8754w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8759w8760w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8765w8766w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8771w8772w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8777w8778w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8783w8784w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8789w8790w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8795w8796w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8801w8802w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8807w8808w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8813w8814w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8819w8820w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8825w8826w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8831w8832w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8837w8838w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8843w8844w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8849w8850w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8855w8856w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8861w8862w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8867w8868w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8873w8874w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8879w8880w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8885w8886w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8891w8892w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8897w8898w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8903w8904w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8909w8910w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8915w8916w
 & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8921w8922w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8927w8928w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8933w8934w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8939w8940w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8945w8946w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8951w8952w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8957w8958w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8963w8964w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8969w8970w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8975w8976w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8981w8982w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8987w8988w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8993w8994w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range8999w9000w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9005w9006w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9011w9012w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9017w9018w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9023w9024w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9029w9030w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9035w9036w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9041w9042w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9047w9048w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9053w9054w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9059w9060w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9065w9066w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9071w9072w & wire_tbl3_taylor_prod_w_lg_w_msb_prod_wo_range9077w9078w);
	result <= ( wire_sum_result(88 DOWNTO 0) & lowest_bits_wo);
	sum_one <= ( wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9975w9976w9977w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9965w9966w9967w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9955w9956w9957w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9945w9946w9947w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9935w9936w9937w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9925w9926w9927w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9915w9916w9917w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9905w9906w9907w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9895w9896w9897w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9885w9886w9887w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9875w9876w9877w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9865w9866w9867w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9855w9856w9857w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9845w9846w9847w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9835w9836w9837w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9825w9826w9827w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9815w9816w9817w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9805w9806w9807w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9795w9796w9797w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9785w9786w9787w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9775w9776w9777w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9765w9766w9767w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9755w9756w9757w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9745w9746w9747w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9735w9736w9737w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9725w9726w9727w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9715w9716w9717w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9705w9706w9707w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9695w9696w9697w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9685w9686w9687w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9675w9676w9677w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9665w9666w9667w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9655w9656w9657w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9645w9646w9647w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9635w9636w9637w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9625w9626w9627w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9615w9616w9617w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9605w9606w9607w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9595w9596w9597w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9585w9586w9587w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9575w9576w9577w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9565w9566w9567w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9555w9556w9557w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9545w9546w9547w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9535w9536w9537w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9525w9526w9527w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9515w9516w9517w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9505w9506w9507w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9495w9496w9497w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9485w9486w9487w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9475w9476w9477w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9465w9466w9467w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9455w9456w9457w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9445w9446w9447w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9435w9436w9437w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9425w9426w9427w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9415w9416w9417w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9405w9406w9407w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9395w9396w9397w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9385w9386w9387w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9375w9376w9377w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9365w9366w9367w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9355w9356w9357w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9345w9346w9347w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9335w9336w9337w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9325w9326w9327w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9315w9316w9317w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9305w9306w9307w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9295w9296w9297w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9285w9286w9287w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9275w9276w9277w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9265w9266w9267w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9255w9256w9257w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9245w9246w9247w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9235w9236w9237w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9225w9226w9227w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9215w9216w9217w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9205w9206w9207w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9195w9196w9197w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9185w9186w9187w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9175w9176w9177w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9165w9166w9167w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9155w9156w9157w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9145w9146w9147w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9135w9136w9137w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9125w9126w9127w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9115w9116w9117w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9105w9106w9107w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9095w9096w9097w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector2_range9083w9084w9085w);
	sum_two <= ( wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10971w10972w10973w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10960w10961w10962w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10949w10950w10951w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10938w10939w10940w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10927w10928w10929w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10916w10917w10918w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10905w10906w10907w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10894w10895w10896w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10883w10884w10885w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10872w10873w10874w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10861w10862w10863w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10850w10851w10852w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10839w10840w10841w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10828w10829w10830w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10817w10818w10819w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10806w10807w10808w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10795w10796w10797w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10784w10785w10786w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10773w10774w10775w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10762w10763w10764w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10751w10752w10753w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10740w10741w10742w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10729w10730w10731w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10718w10719w10720w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10707w10708w10709w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10696w10697w10698w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10685w10686w10687w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10674w10675w10676w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10663w10664w10665w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10652w10653w10654w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10641w10642w10643w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10630w10631w10632w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10619w10620w10621w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10608w10609w10610w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10597w10598w10599w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10586w10587w10588w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10575w10576w10577w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10564w10565w10566w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10553w10554w10555w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10542w10543w10544w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10531w10532w10533w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10520w10521w10522w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10509w10510w10511w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10498w10499w10500w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10487w10488w10489w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10476w10477w10478w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10465w10466w10467w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10454w10455w10456w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10443w10444w10445w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10432w10433w10434w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10421w10422w10423w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10410w10411w10412w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10399w10400w10401w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10388w10389w10390w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10377w10378w10379w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10366w10367w10368w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10355w10356w10357w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10344w10345w10346w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10333w10334w10335w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10322w10323w10324w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10311w10312w10313w
 & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10300w10301w10302w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10289w10290w10291w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10278w10279w10280w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10267w10268w10269w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10256w10257w10258w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10245w10246w10247w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10234w10235w10236w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10223w10224w10225w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10212w10213w10214w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10201w10202w10203w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10190w10191w10192w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10179w10180w10181w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10168w10169w10170w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10157w10158w10159w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10146w10147w10148w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10135w10136w10137w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10124w10125w10126w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10113w10114w10115w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10102w10103w10104w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10091w10092w10093w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10080w10081w10082w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10069w10070w10071w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10058w10059w10060w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10047w10048w10049w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10036w10037w10038w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10025w10026w10027w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10014w10015w10016w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range10003w10004w10005w & wire_tbl3_taylor_prod_w_lg_w_lg_w_vector1_range9990w9991w9992w);
	sum_two_wo <= sum_two_reg0;
	vector1 <= ( msb_prod_wo & lsb_prod_wo(61 DOWNTO 31));
	vector2 <= ( "00000000000000000000000000" & mid_prod_wo);
	wire_a <= dataa;
	wire_b <= datab;
	wire_tbl3_taylor_prod_w_car_one_adj_range9988w(0) <= car_one_adj(0);
	wire_tbl3_taylor_prod_w_car_one_adj_range10101w(0) <= car_one_adj(10);
	wire_tbl3_taylor_prod_w_car_one_adj_range10112w(0) <= car_one_adj(11);
	wire_tbl3_taylor_prod_w_car_one_adj_range10123w(0) <= car_one_adj(12);
	wire_tbl3_taylor_prod_w_car_one_adj_range10134w(0) <= car_one_adj(13);
	wire_tbl3_taylor_prod_w_car_one_adj_range10145w(0) <= car_one_adj(14);
	wire_tbl3_taylor_prod_w_car_one_adj_range10156w(0) <= car_one_adj(15);
	wire_tbl3_taylor_prod_w_car_one_adj_range10167w(0) <= car_one_adj(16);
	wire_tbl3_taylor_prod_w_car_one_adj_range10178w(0) <= car_one_adj(17);
	wire_tbl3_taylor_prod_w_car_one_adj_range10189w(0) <= car_one_adj(18);
	wire_tbl3_taylor_prod_w_car_one_adj_range10200w(0) <= car_one_adj(19);
	wire_tbl3_taylor_prod_w_car_one_adj_range10002w(0) <= car_one_adj(1);
	wire_tbl3_taylor_prod_w_car_one_adj_range10211w(0) <= car_one_adj(20);
	wire_tbl3_taylor_prod_w_car_one_adj_range10222w(0) <= car_one_adj(21);
	wire_tbl3_taylor_prod_w_car_one_adj_range10233w(0) <= car_one_adj(22);
	wire_tbl3_taylor_prod_w_car_one_adj_range10244w(0) <= car_one_adj(23);
	wire_tbl3_taylor_prod_w_car_one_adj_range10255w(0) <= car_one_adj(24);
	wire_tbl3_taylor_prod_w_car_one_adj_range10266w(0) <= car_one_adj(25);
	wire_tbl3_taylor_prod_w_car_one_adj_range10277w(0) <= car_one_adj(26);
	wire_tbl3_taylor_prod_w_car_one_adj_range10288w(0) <= car_one_adj(27);
	wire_tbl3_taylor_prod_w_car_one_adj_range10299w(0) <= car_one_adj(28);
	wire_tbl3_taylor_prod_w_car_one_adj_range10310w(0) <= car_one_adj(29);
	wire_tbl3_taylor_prod_w_car_one_adj_range10013w(0) <= car_one_adj(2);
	wire_tbl3_taylor_prod_w_car_one_adj_range10321w(0) <= car_one_adj(30);
	wire_tbl3_taylor_prod_w_car_one_adj_range10332w(0) <= car_one_adj(31);
	wire_tbl3_taylor_prod_w_car_one_adj_range10343w(0) <= car_one_adj(32);
	wire_tbl3_taylor_prod_w_car_one_adj_range10354w(0) <= car_one_adj(33);
	wire_tbl3_taylor_prod_w_car_one_adj_range10365w(0) <= car_one_adj(34);
	wire_tbl3_taylor_prod_w_car_one_adj_range10376w(0) <= car_one_adj(35);
	wire_tbl3_taylor_prod_w_car_one_adj_range10387w(0) <= car_one_adj(36);
	wire_tbl3_taylor_prod_w_car_one_adj_range10398w(0) <= car_one_adj(37);
	wire_tbl3_taylor_prod_w_car_one_adj_range10409w(0) <= car_one_adj(38);
	wire_tbl3_taylor_prod_w_car_one_adj_range10420w(0) <= car_one_adj(39);
	wire_tbl3_taylor_prod_w_car_one_adj_range10024w(0) <= car_one_adj(3);
	wire_tbl3_taylor_prod_w_car_one_adj_range10431w(0) <= car_one_adj(40);
	wire_tbl3_taylor_prod_w_car_one_adj_range10442w(0) <= car_one_adj(41);
	wire_tbl3_taylor_prod_w_car_one_adj_range10453w(0) <= car_one_adj(42);
	wire_tbl3_taylor_prod_w_car_one_adj_range10464w(0) <= car_one_adj(43);
	wire_tbl3_taylor_prod_w_car_one_adj_range10475w(0) <= car_one_adj(44);
	wire_tbl3_taylor_prod_w_car_one_adj_range10486w(0) <= car_one_adj(45);
	wire_tbl3_taylor_prod_w_car_one_adj_range10497w(0) <= car_one_adj(46);
	wire_tbl3_taylor_prod_w_car_one_adj_range10508w(0) <= car_one_adj(47);
	wire_tbl3_taylor_prod_w_car_one_adj_range10519w(0) <= car_one_adj(48);
	wire_tbl3_taylor_prod_w_car_one_adj_range10530w(0) <= car_one_adj(49);
	wire_tbl3_taylor_prod_w_car_one_adj_range10035w(0) <= car_one_adj(4);
	wire_tbl3_taylor_prod_w_car_one_adj_range10541w(0) <= car_one_adj(50);
	wire_tbl3_taylor_prod_w_car_one_adj_range10552w(0) <= car_one_adj(51);
	wire_tbl3_taylor_prod_w_car_one_adj_range10563w(0) <= car_one_adj(52);
	wire_tbl3_taylor_prod_w_car_one_adj_range10574w(0) <= car_one_adj(53);
	wire_tbl3_taylor_prod_w_car_one_adj_range10585w(0) <= car_one_adj(54);
	wire_tbl3_taylor_prod_w_car_one_adj_range10596w(0) <= car_one_adj(55);
	wire_tbl3_taylor_prod_w_car_one_adj_range10607w(0) <= car_one_adj(56);
	wire_tbl3_taylor_prod_w_car_one_adj_range10618w(0) <= car_one_adj(57);
	wire_tbl3_taylor_prod_w_car_one_adj_range10629w(0) <= car_one_adj(58);
	wire_tbl3_taylor_prod_w_car_one_adj_range10640w(0) <= car_one_adj(59);
	wire_tbl3_taylor_prod_w_car_one_adj_range10046w(0) <= car_one_adj(5);
	wire_tbl3_taylor_prod_w_car_one_adj_range10651w(0) <= car_one_adj(60);
	wire_tbl3_taylor_prod_w_car_one_adj_range10662w(0) <= car_one_adj(61);
	wire_tbl3_taylor_prod_w_car_one_adj_range10673w(0) <= car_one_adj(62);
	wire_tbl3_taylor_prod_w_car_one_adj_range10684w(0) <= car_one_adj(63);
	wire_tbl3_taylor_prod_w_car_one_adj_range10695w(0) <= car_one_adj(64);
	wire_tbl3_taylor_prod_w_car_one_adj_range10706w(0) <= car_one_adj(65);
	wire_tbl3_taylor_prod_w_car_one_adj_range10717w(0) <= car_one_adj(66);
	wire_tbl3_taylor_prod_w_car_one_adj_range10728w(0) <= car_one_adj(67);
	wire_tbl3_taylor_prod_w_car_one_adj_range10739w(0) <= car_one_adj(68);
	wire_tbl3_taylor_prod_w_car_one_adj_range10750w(0) <= car_one_adj(69);
	wire_tbl3_taylor_prod_w_car_one_adj_range10057w(0) <= car_one_adj(6);
	wire_tbl3_taylor_prod_w_car_one_adj_range10761w(0) <= car_one_adj(70);
	wire_tbl3_taylor_prod_w_car_one_adj_range10772w(0) <= car_one_adj(71);
	wire_tbl3_taylor_prod_w_car_one_adj_range10783w(0) <= car_one_adj(72);
	wire_tbl3_taylor_prod_w_car_one_adj_range10794w(0) <= car_one_adj(73);
	wire_tbl3_taylor_prod_w_car_one_adj_range10805w(0) <= car_one_adj(74);
	wire_tbl3_taylor_prod_w_car_one_adj_range10816w(0) <= car_one_adj(75);
	wire_tbl3_taylor_prod_w_car_one_adj_range10827w(0) <= car_one_adj(76);
	wire_tbl3_taylor_prod_w_car_one_adj_range10838w(0) <= car_one_adj(77);
	wire_tbl3_taylor_prod_w_car_one_adj_range10849w(0) <= car_one_adj(78);
	wire_tbl3_taylor_prod_w_car_one_adj_range10860w(0) <= car_one_adj(79);
	wire_tbl3_taylor_prod_w_car_one_adj_range10068w(0) <= car_one_adj(7);
	wire_tbl3_taylor_prod_w_car_one_adj_range10871w(0) <= car_one_adj(80);
	wire_tbl3_taylor_prod_w_car_one_adj_range10882w(0) <= car_one_adj(81);
	wire_tbl3_taylor_prod_w_car_one_adj_range10893w(0) <= car_one_adj(82);
	wire_tbl3_taylor_prod_w_car_one_adj_range10904w(0) <= car_one_adj(83);
	wire_tbl3_taylor_prod_w_car_one_adj_range10915w(0) <= car_one_adj(84);
	wire_tbl3_taylor_prod_w_car_one_adj_range10926w(0) <= car_one_adj(85);
	wire_tbl3_taylor_prod_w_car_one_adj_range10937w(0) <= car_one_adj(86);
	wire_tbl3_taylor_prod_w_car_one_adj_range10948w(0) <= car_one_adj(87);
	wire_tbl3_taylor_prod_w_car_one_adj_range10959w(0) <= car_one_adj(88);
	wire_tbl3_taylor_prod_w_car_one_adj_range10970w(0) <= car_one_adj(89);
	wire_tbl3_taylor_prod_w_car_one_adj_range10079w(0) <= car_one_adj(8);
	wire_tbl3_taylor_prod_w_car_one_adj_range10090w(0) <= car_one_adj(9);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9080w(0) <= lsb_prod_wo(0);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9020w(0) <= lsb_prod_wo(10);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9014w(0) <= lsb_prod_wo(11);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9008w(0) <= lsb_prod_wo(12);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9002w(0) <= lsb_prod_wo(13);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8996w(0) <= lsb_prod_wo(14);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8990w(0) <= lsb_prod_wo(15);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8984w(0) <= lsb_prod_wo(16);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8978w(0) <= lsb_prod_wo(17);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8972w(0) <= lsb_prod_wo(18);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8966w(0) <= lsb_prod_wo(19);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9074w(0) <= lsb_prod_wo(1);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8960w(0) <= lsb_prod_wo(20);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8954w(0) <= lsb_prod_wo(21);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8948w(0) <= lsb_prod_wo(22);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8942w(0) <= lsb_prod_wo(23);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8936w(0) <= lsb_prod_wo(24);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8930w(0) <= lsb_prod_wo(25);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8924w(0) <= lsb_prod_wo(26);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8918w(0) <= lsb_prod_wo(27);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8912w(0) <= lsb_prod_wo(28);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8906w(0) <= lsb_prod_wo(29);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9068w(0) <= lsb_prod_wo(2);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8900w(0) <= lsb_prod_wo(30);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8894w(0) <= lsb_prod_wo(31);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8888w(0) <= lsb_prod_wo(32);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8882w(0) <= lsb_prod_wo(33);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8876w(0) <= lsb_prod_wo(34);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8870w(0) <= lsb_prod_wo(35);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8864w(0) <= lsb_prod_wo(36);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8858w(0) <= lsb_prod_wo(37);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8852w(0) <= lsb_prod_wo(38);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8846w(0) <= lsb_prod_wo(39);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9062w(0) <= lsb_prod_wo(3);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8840w(0) <= lsb_prod_wo(40);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8834w(0) <= lsb_prod_wo(41);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8828w(0) <= lsb_prod_wo(42);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8822w(0) <= lsb_prod_wo(43);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8816w(0) <= lsb_prod_wo(44);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8810w(0) <= lsb_prod_wo(45);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8804w(0) <= lsb_prod_wo(46);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8798w(0) <= lsb_prod_wo(47);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8792w(0) <= lsb_prod_wo(48);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8786w(0) <= lsb_prod_wo(49);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9056w(0) <= lsb_prod_wo(4);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8780w(0) <= lsb_prod_wo(50);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8774w(0) <= lsb_prod_wo(51);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8768w(0) <= lsb_prod_wo(52);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8762w(0) <= lsb_prod_wo(53);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8756w(0) <= lsb_prod_wo(54);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8750w(0) <= lsb_prod_wo(55);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8744w(0) <= lsb_prod_wo(56);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8738w(0) <= lsb_prod_wo(57);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8732w(0) <= lsb_prod_wo(58);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8726w(0) <= lsb_prod_wo(59);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9050w(0) <= lsb_prod_wo(5);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8721w(0) <= lsb_prod_wo(60);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range8716w(0) <= lsb_prod_wo(61);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9044w(0) <= lsb_prod_wo(6);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9038w(0) <= lsb_prod_wo(7);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9032w(0) <= lsb_prod_wo(8);
	wire_tbl3_taylor_prod_w_lsb_prod_wo_range9026w(0) <= lsb_prod_wo(9);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9077w(0) <= msb_prod_wo(0);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9017w(0) <= msb_prod_wo(10);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9011w(0) <= msb_prod_wo(11);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9005w(0) <= msb_prod_wo(12);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8999w(0) <= msb_prod_wo(13);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8993w(0) <= msb_prod_wo(14);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8987w(0) <= msb_prod_wo(15);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8981w(0) <= msb_prod_wo(16);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8975w(0) <= msb_prod_wo(17);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8969w(0) <= msb_prod_wo(18);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8963w(0) <= msb_prod_wo(19);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9071w(0) <= msb_prod_wo(1);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8957w(0) <= msb_prod_wo(20);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8951w(0) <= msb_prod_wo(21);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8945w(0) <= msb_prod_wo(22);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8939w(0) <= msb_prod_wo(23);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8933w(0) <= msb_prod_wo(24);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8927w(0) <= msb_prod_wo(25);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8921w(0) <= msb_prod_wo(26);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8915w(0) <= msb_prod_wo(27);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8909w(0) <= msb_prod_wo(28);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8903w(0) <= msb_prod_wo(29);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9065w(0) <= msb_prod_wo(2);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8897w(0) <= msb_prod_wo(30);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8891w(0) <= msb_prod_wo(31);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8885w(0) <= msb_prod_wo(32);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8879w(0) <= msb_prod_wo(33);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8873w(0) <= msb_prod_wo(34);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8867w(0) <= msb_prod_wo(35);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8861w(0) <= msb_prod_wo(36);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8855w(0) <= msb_prod_wo(37);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8849w(0) <= msb_prod_wo(38);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8843w(0) <= msb_prod_wo(39);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9059w(0) <= msb_prod_wo(3);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8837w(0) <= msb_prod_wo(40);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8831w(0) <= msb_prod_wo(41);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8825w(0) <= msb_prod_wo(42);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8819w(0) <= msb_prod_wo(43);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8813w(0) <= msb_prod_wo(44);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8807w(0) <= msb_prod_wo(45);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8801w(0) <= msb_prod_wo(46);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8795w(0) <= msb_prod_wo(47);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8789w(0) <= msb_prod_wo(48);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8783w(0) <= msb_prod_wo(49);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9053w(0) <= msb_prod_wo(4);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8777w(0) <= msb_prod_wo(50);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8771w(0) <= msb_prod_wo(51);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8765w(0) <= msb_prod_wo(52);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8759w(0) <= msb_prod_wo(53);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8753w(0) <= msb_prod_wo(54);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8747w(0) <= msb_prod_wo(55);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8741w(0) <= msb_prod_wo(56);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8735w(0) <= msb_prod_wo(57);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range8729w(0) <= msb_prod_wo(58);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9047w(0) <= msb_prod_wo(5);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9041w(0) <= msb_prod_wo(6);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9035w(0) <= msb_prod_wo(7);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9029w(0) <= msb_prod_wo(8);
	wire_tbl3_taylor_prod_w_msb_prod_wo_range9023w(0) <= msb_prod_wo(9);
	wire_tbl3_taylor_prod_w_neg_lsb_range9082w(0) <= neg_lsb(0);
	wire_tbl3_taylor_prod_w_neg_lsb_range9022w(0) <= neg_lsb(10);
	wire_tbl3_taylor_prod_w_neg_lsb_range9016w(0) <= neg_lsb(11);
	wire_tbl3_taylor_prod_w_neg_lsb_range9010w(0) <= neg_lsb(12);
	wire_tbl3_taylor_prod_w_neg_lsb_range9004w(0) <= neg_lsb(13);
	wire_tbl3_taylor_prod_w_neg_lsb_range8998w(0) <= neg_lsb(14);
	wire_tbl3_taylor_prod_w_neg_lsb_range8992w(0) <= neg_lsb(15);
	wire_tbl3_taylor_prod_w_neg_lsb_range8986w(0) <= neg_lsb(16);
	wire_tbl3_taylor_prod_w_neg_lsb_range8980w(0) <= neg_lsb(17);
	wire_tbl3_taylor_prod_w_neg_lsb_range8974w(0) <= neg_lsb(18);
	wire_tbl3_taylor_prod_w_neg_lsb_range8968w(0) <= neg_lsb(19);
	wire_tbl3_taylor_prod_w_neg_lsb_range9076w(0) <= neg_lsb(1);
	wire_tbl3_taylor_prod_w_neg_lsb_range8962w(0) <= neg_lsb(20);
	wire_tbl3_taylor_prod_w_neg_lsb_range8956w(0) <= neg_lsb(21);
	wire_tbl3_taylor_prod_w_neg_lsb_range8950w(0) <= neg_lsb(22);
	wire_tbl3_taylor_prod_w_neg_lsb_range8944w(0) <= neg_lsb(23);
	wire_tbl3_taylor_prod_w_neg_lsb_range8938w(0) <= neg_lsb(24);
	wire_tbl3_taylor_prod_w_neg_lsb_range8932w(0) <= neg_lsb(25);
	wire_tbl3_taylor_prod_w_neg_lsb_range8926w(0) <= neg_lsb(26);
	wire_tbl3_taylor_prod_w_neg_lsb_range8920w(0) <= neg_lsb(27);
	wire_tbl3_taylor_prod_w_neg_lsb_range8914w(0) <= neg_lsb(28);
	wire_tbl3_taylor_prod_w_neg_lsb_range8908w(0) <= neg_lsb(29);
	wire_tbl3_taylor_prod_w_neg_lsb_range9070w(0) <= neg_lsb(2);
	wire_tbl3_taylor_prod_w_neg_lsb_range8902w(0) <= neg_lsb(30);
	wire_tbl3_taylor_prod_w_neg_lsb_range8896w(0) <= neg_lsb(31);
	wire_tbl3_taylor_prod_w_neg_lsb_range8890w(0) <= neg_lsb(32);
	wire_tbl3_taylor_prod_w_neg_lsb_range8884w(0) <= neg_lsb(33);
	wire_tbl3_taylor_prod_w_neg_lsb_range8878w(0) <= neg_lsb(34);
	wire_tbl3_taylor_prod_w_neg_lsb_range8872w(0) <= neg_lsb(35);
	wire_tbl3_taylor_prod_w_neg_lsb_range8866w(0) <= neg_lsb(36);
	wire_tbl3_taylor_prod_w_neg_lsb_range8860w(0) <= neg_lsb(37);
	wire_tbl3_taylor_prod_w_neg_lsb_range8854w(0) <= neg_lsb(38);
	wire_tbl3_taylor_prod_w_neg_lsb_range8848w(0) <= neg_lsb(39);
	wire_tbl3_taylor_prod_w_neg_lsb_range9064w(0) <= neg_lsb(3);
	wire_tbl3_taylor_prod_w_neg_lsb_range8842w(0) <= neg_lsb(40);
	wire_tbl3_taylor_prod_w_neg_lsb_range8836w(0) <= neg_lsb(41);
	wire_tbl3_taylor_prod_w_neg_lsb_range8830w(0) <= neg_lsb(42);
	wire_tbl3_taylor_prod_w_neg_lsb_range8824w(0) <= neg_lsb(43);
	wire_tbl3_taylor_prod_w_neg_lsb_range8818w(0) <= neg_lsb(44);
	wire_tbl3_taylor_prod_w_neg_lsb_range8812w(0) <= neg_lsb(45);
	wire_tbl3_taylor_prod_w_neg_lsb_range8806w(0) <= neg_lsb(46);
	wire_tbl3_taylor_prod_w_neg_lsb_range8800w(0) <= neg_lsb(47);
	wire_tbl3_taylor_prod_w_neg_lsb_range8794w(0) <= neg_lsb(48);
	wire_tbl3_taylor_prod_w_neg_lsb_range8788w(0) <= neg_lsb(49);
	wire_tbl3_taylor_prod_w_neg_lsb_range9058w(0) <= neg_lsb(4);
	wire_tbl3_taylor_prod_w_neg_lsb_range8782w(0) <= neg_lsb(50);
	wire_tbl3_taylor_prod_w_neg_lsb_range8776w(0) <= neg_lsb(51);
	wire_tbl3_taylor_prod_w_neg_lsb_range8770w(0) <= neg_lsb(52);
	wire_tbl3_taylor_prod_w_neg_lsb_range8764w(0) <= neg_lsb(53);
	wire_tbl3_taylor_prod_w_neg_lsb_range8758w(0) <= neg_lsb(54);
	wire_tbl3_taylor_prod_w_neg_lsb_range8752w(0) <= neg_lsb(55);
	wire_tbl3_taylor_prod_w_neg_lsb_range8746w(0) <= neg_lsb(56);
	wire_tbl3_taylor_prod_w_neg_lsb_range8740w(0) <= neg_lsb(57);
	wire_tbl3_taylor_prod_w_neg_lsb_range8734w(0) <= neg_lsb(58);
	wire_tbl3_taylor_prod_w_neg_lsb_range8728w(0) <= neg_lsb(59);
	wire_tbl3_taylor_prod_w_neg_lsb_range9052w(0) <= neg_lsb(5);
	wire_tbl3_taylor_prod_w_neg_lsb_range8723w(0) <= neg_lsb(60);
	wire_tbl3_taylor_prod_w_neg_lsb_range8718w(0) <= neg_lsb(61);
	wire_tbl3_taylor_prod_w_neg_lsb_range8712w(0) <= neg_lsb(62);
	wire_tbl3_taylor_prod_w_neg_lsb_range8708w(0) <= neg_lsb(63);
	wire_tbl3_taylor_prod_w_neg_lsb_range8704w(0) <= neg_lsb(64);
	wire_tbl3_taylor_prod_w_neg_lsb_range8700w(0) <= neg_lsb(65);
	wire_tbl3_taylor_prod_w_neg_lsb_range8696w(0) <= neg_lsb(66);
	wire_tbl3_taylor_prod_w_neg_lsb_range8692w(0) <= neg_lsb(67);
	wire_tbl3_taylor_prod_w_neg_lsb_range8688w(0) <= neg_lsb(68);
	wire_tbl3_taylor_prod_w_neg_lsb_range8684w(0) <= neg_lsb(69);
	wire_tbl3_taylor_prod_w_neg_lsb_range9046w(0) <= neg_lsb(6);
	wire_tbl3_taylor_prod_w_neg_lsb_range8680w(0) <= neg_lsb(70);
	wire_tbl3_taylor_prod_w_neg_lsb_range8676w(0) <= neg_lsb(71);
	wire_tbl3_taylor_prod_w_neg_lsb_range8672w(0) <= neg_lsb(72);
	wire_tbl3_taylor_prod_w_neg_lsb_range8668w(0) <= neg_lsb(73);
	wire_tbl3_taylor_prod_w_neg_lsb_range8664w(0) <= neg_lsb(74);
	wire_tbl3_taylor_prod_w_neg_lsb_range8660w(0) <= neg_lsb(75);
	wire_tbl3_taylor_prod_w_neg_lsb_range8656w(0) <= neg_lsb(76);
	wire_tbl3_taylor_prod_w_neg_lsb_range8652w(0) <= neg_lsb(77);
	wire_tbl3_taylor_prod_w_neg_lsb_range8648w(0) <= neg_lsb(78);
	wire_tbl3_taylor_prod_w_neg_lsb_range8644w(0) <= neg_lsb(79);
	wire_tbl3_taylor_prod_w_neg_lsb_range9040w(0) <= neg_lsb(7);
	wire_tbl3_taylor_prod_w_neg_lsb_range8640w(0) <= neg_lsb(80);
	wire_tbl3_taylor_prod_w_neg_lsb_range8636w(0) <= neg_lsb(81);
	wire_tbl3_taylor_prod_w_neg_lsb_range8632w(0) <= neg_lsb(82);
	wire_tbl3_taylor_prod_w_neg_lsb_range8628w(0) <= neg_lsb(83);
	wire_tbl3_taylor_prod_w_neg_lsb_range8624w(0) <= neg_lsb(84);
	wire_tbl3_taylor_prod_w_neg_lsb_range8620w(0) <= neg_lsb(85);
	wire_tbl3_taylor_prod_w_neg_lsb_range8616w(0) <= neg_lsb(86);
	wire_tbl3_taylor_prod_w_neg_lsb_range8612w(0) <= neg_lsb(87);
	wire_tbl3_taylor_prod_w_neg_lsb_range8608w(0) <= neg_lsb(88);
	wire_tbl3_taylor_prod_w_neg_lsb_range8603w(0) <= neg_lsb(89);
	wire_tbl3_taylor_prod_w_neg_lsb_range9034w(0) <= neg_lsb(8);
	wire_tbl3_taylor_prod_w_neg_lsb_range9028w(0) <= neg_lsb(9);
	wire_tbl3_taylor_prod_w_neg_msb_range9079w(0) <= neg_msb(0);
	wire_tbl3_taylor_prod_w_neg_msb_range9019w(0) <= neg_msb(10);
	wire_tbl3_taylor_prod_w_neg_msb_range9013w(0) <= neg_msb(11);
	wire_tbl3_taylor_prod_w_neg_msb_range9007w(0) <= neg_msb(12);
	wire_tbl3_taylor_prod_w_neg_msb_range9001w(0) <= neg_msb(13);
	wire_tbl3_taylor_prod_w_neg_msb_range8995w(0) <= neg_msb(14);
	wire_tbl3_taylor_prod_w_neg_msb_range8989w(0) <= neg_msb(15);
	wire_tbl3_taylor_prod_w_neg_msb_range8983w(0) <= neg_msb(16);
	wire_tbl3_taylor_prod_w_neg_msb_range8977w(0) <= neg_msb(17);
	wire_tbl3_taylor_prod_w_neg_msb_range8971w(0) <= neg_msb(18);
	wire_tbl3_taylor_prod_w_neg_msb_range8965w(0) <= neg_msb(19);
	wire_tbl3_taylor_prod_w_neg_msb_range9073w(0) <= neg_msb(1);
	wire_tbl3_taylor_prod_w_neg_msb_range8959w(0) <= neg_msb(20);
	wire_tbl3_taylor_prod_w_neg_msb_range8953w(0) <= neg_msb(21);
	wire_tbl3_taylor_prod_w_neg_msb_range8947w(0) <= neg_msb(22);
	wire_tbl3_taylor_prod_w_neg_msb_range8941w(0) <= neg_msb(23);
	wire_tbl3_taylor_prod_w_neg_msb_range8935w(0) <= neg_msb(24);
	wire_tbl3_taylor_prod_w_neg_msb_range8929w(0) <= neg_msb(25);
	wire_tbl3_taylor_prod_w_neg_msb_range8923w(0) <= neg_msb(26);
	wire_tbl3_taylor_prod_w_neg_msb_range8917w(0) <= neg_msb(27);
	wire_tbl3_taylor_prod_w_neg_msb_range8911w(0) <= neg_msb(28);
	wire_tbl3_taylor_prod_w_neg_msb_range8905w(0) <= neg_msb(29);
	wire_tbl3_taylor_prod_w_neg_msb_range9067w(0) <= neg_msb(2);
	wire_tbl3_taylor_prod_w_neg_msb_range8899w(0) <= neg_msb(30);
	wire_tbl3_taylor_prod_w_neg_msb_range8893w(0) <= neg_msb(31);
	wire_tbl3_taylor_prod_w_neg_msb_range8887w(0) <= neg_msb(32);
	wire_tbl3_taylor_prod_w_neg_msb_range8881w(0) <= neg_msb(33);
	wire_tbl3_taylor_prod_w_neg_msb_range8875w(0) <= neg_msb(34);
	wire_tbl3_taylor_prod_w_neg_msb_range8869w(0) <= neg_msb(35);
	wire_tbl3_taylor_prod_w_neg_msb_range8863w(0) <= neg_msb(36);
	wire_tbl3_taylor_prod_w_neg_msb_range8857w(0) <= neg_msb(37);
	wire_tbl3_taylor_prod_w_neg_msb_range8851w(0) <= neg_msb(38);
	wire_tbl3_taylor_prod_w_neg_msb_range8845w(0) <= neg_msb(39);
	wire_tbl3_taylor_prod_w_neg_msb_range9061w(0) <= neg_msb(3);
	wire_tbl3_taylor_prod_w_neg_msb_range8839w(0) <= neg_msb(40);
	wire_tbl3_taylor_prod_w_neg_msb_range8833w(0) <= neg_msb(41);
	wire_tbl3_taylor_prod_w_neg_msb_range8827w(0) <= neg_msb(42);
	wire_tbl3_taylor_prod_w_neg_msb_range8821w(0) <= neg_msb(43);
	wire_tbl3_taylor_prod_w_neg_msb_range8815w(0) <= neg_msb(44);
	wire_tbl3_taylor_prod_w_neg_msb_range8809w(0) <= neg_msb(45);
	wire_tbl3_taylor_prod_w_neg_msb_range8803w(0) <= neg_msb(46);
	wire_tbl3_taylor_prod_w_neg_msb_range8797w(0) <= neg_msb(47);
	wire_tbl3_taylor_prod_w_neg_msb_range8791w(0) <= neg_msb(48);
	wire_tbl3_taylor_prod_w_neg_msb_range8785w(0) <= neg_msb(49);
	wire_tbl3_taylor_prod_w_neg_msb_range9055w(0) <= neg_msb(4);
	wire_tbl3_taylor_prod_w_neg_msb_range8779w(0) <= neg_msb(50);
	wire_tbl3_taylor_prod_w_neg_msb_range8773w(0) <= neg_msb(51);
	wire_tbl3_taylor_prod_w_neg_msb_range8767w(0) <= neg_msb(52);
	wire_tbl3_taylor_prod_w_neg_msb_range8761w(0) <= neg_msb(53);
	wire_tbl3_taylor_prod_w_neg_msb_range8755w(0) <= neg_msb(54);
	wire_tbl3_taylor_prod_w_neg_msb_range8749w(0) <= neg_msb(55);
	wire_tbl3_taylor_prod_w_neg_msb_range8743w(0) <= neg_msb(56);
	wire_tbl3_taylor_prod_w_neg_msb_range8737w(0) <= neg_msb(57);
	wire_tbl3_taylor_prod_w_neg_msb_range8731w(0) <= neg_msb(58);
	wire_tbl3_taylor_prod_w_neg_msb_range8724w(0) <= neg_msb(59);
	wire_tbl3_taylor_prod_w_neg_msb_range9049w(0) <= neg_msb(5);
	wire_tbl3_taylor_prod_w_neg_msb_range8719w(0) <= neg_msb(60);
	wire_tbl3_taylor_prod_w_neg_msb_range8714w(0) <= neg_msb(61);
	wire_tbl3_taylor_prod_w_neg_msb_range8710w(0) <= neg_msb(62);
	wire_tbl3_taylor_prod_w_neg_msb_range8706w(0) <= neg_msb(63);
	wire_tbl3_taylor_prod_w_neg_msb_range8702w(0) <= neg_msb(64);
	wire_tbl3_taylor_prod_w_neg_msb_range8698w(0) <= neg_msb(65);
	wire_tbl3_taylor_prod_w_neg_msb_range8694w(0) <= neg_msb(66);
	wire_tbl3_taylor_prod_w_neg_msb_range8690w(0) <= neg_msb(67);
	wire_tbl3_taylor_prod_w_neg_msb_range8686w(0) <= neg_msb(68);
	wire_tbl3_taylor_prod_w_neg_msb_range8682w(0) <= neg_msb(69);
	wire_tbl3_taylor_prod_w_neg_msb_range9043w(0) <= neg_msb(6);
	wire_tbl3_taylor_prod_w_neg_msb_range8678w(0) <= neg_msb(70);
	wire_tbl3_taylor_prod_w_neg_msb_range8674w(0) <= neg_msb(71);
	wire_tbl3_taylor_prod_w_neg_msb_range8670w(0) <= neg_msb(72);
	wire_tbl3_taylor_prod_w_neg_msb_range8666w(0) <= neg_msb(73);
	wire_tbl3_taylor_prod_w_neg_msb_range8662w(0) <= neg_msb(74);
	wire_tbl3_taylor_prod_w_neg_msb_range8658w(0) <= neg_msb(75);
	wire_tbl3_taylor_prod_w_neg_msb_range8654w(0) <= neg_msb(76);
	wire_tbl3_taylor_prod_w_neg_msb_range8650w(0) <= neg_msb(77);
	wire_tbl3_taylor_prod_w_neg_msb_range8646w(0) <= neg_msb(78);
	wire_tbl3_taylor_prod_w_neg_msb_range8642w(0) <= neg_msb(79);
	wire_tbl3_taylor_prod_w_neg_msb_range9037w(0) <= neg_msb(7);
	wire_tbl3_taylor_prod_w_neg_msb_range8638w(0) <= neg_msb(80);
	wire_tbl3_taylor_prod_w_neg_msb_range8634w(0) <= neg_msb(81);
	wire_tbl3_taylor_prod_w_neg_msb_range8630w(0) <= neg_msb(82);
	wire_tbl3_taylor_prod_w_neg_msb_range8626w(0) <= neg_msb(83);
	wire_tbl3_taylor_prod_w_neg_msb_range8622w(0) <= neg_msb(84);
	wire_tbl3_taylor_prod_w_neg_msb_range8618w(0) <= neg_msb(85);
	wire_tbl3_taylor_prod_w_neg_msb_range8614w(0) <= neg_msb(86);
	wire_tbl3_taylor_prod_w_neg_msb_range8610w(0) <= neg_msb(87);
	wire_tbl3_taylor_prod_w_neg_msb_range8606w(0) <= neg_msb(88);
	wire_tbl3_taylor_prod_w_neg_msb_range8600w(0) <= neg_msb(89);
	wire_tbl3_taylor_prod_w_neg_msb_range9031w(0) <= neg_msb(8);
	wire_tbl3_taylor_prod_w_neg_msb_range9025w(0) <= neg_msb(9);
	wire_tbl3_taylor_prod_w_sum_one_range9086w(0) <= sum_one(0);
	wire_tbl3_taylor_prod_w_sum_one_range9188w(0) <= sum_one(10);
	wire_tbl3_taylor_prod_w_sum_one_range9198w(0) <= sum_one(11);
	wire_tbl3_taylor_prod_w_sum_one_range9208w(0) <= sum_one(12);
	wire_tbl3_taylor_prod_w_sum_one_range9218w(0) <= sum_one(13);
	wire_tbl3_taylor_prod_w_sum_one_range9228w(0) <= sum_one(14);
	wire_tbl3_taylor_prod_w_sum_one_range9238w(0) <= sum_one(15);
	wire_tbl3_taylor_prod_w_sum_one_range9248w(0) <= sum_one(16);
	wire_tbl3_taylor_prod_w_sum_one_range9258w(0) <= sum_one(17);
	wire_tbl3_taylor_prod_w_sum_one_range9268w(0) <= sum_one(18);
	wire_tbl3_taylor_prod_w_sum_one_range9278w(0) <= sum_one(19);
	wire_tbl3_taylor_prod_w_sum_one_range9098w(0) <= sum_one(1);
	wire_tbl3_taylor_prod_w_sum_one_range9288w(0) <= sum_one(20);
	wire_tbl3_taylor_prod_w_sum_one_range9298w(0) <= sum_one(21);
	wire_tbl3_taylor_prod_w_sum_one_range9308w(0) <= sum_one(22);
	wire_tbl3_taylor_prod_w_sum_one_range9318w(0) <= sum_one(23);
	wire_tbl3_taylor_prod_w_sum_one_range9328w(0) <= sum_one(24);
	wire_tbl3_taylor_prod_w_sum_one_range9338w(0) <= sum_one(25);
	wire_tbl3_taylor_prod_w_sum_one_range9348w(0) <= sum_one(26);
	wire_tbl3_taylor_prod_w_sum_one_range9358w(0) <= sum_one(27);
	wire_tbl3_taylor_prod_w_sum_one_range9368w(0) <= sum_one(28);
	wire_tbl3_taylor_prod_w_sum_one_range9378w(0) <= sum_one(29);
	wire_tbl3_taylor_prod_w_sum_one_range9108w(0) <= sum_one(2);
	wire_tbl3_taylor_prod_w_sum_one_range9388w(0) <= sum_one(30);
	wire_tbl3_taylor_prod_w_sum_one_range9398w(0) <= sum_one(31);
	wire_tbl3_taylor_prod_w_sum_one_range9408w(0) <= sum_one(32);
	wire_tbl3_taylor_prod_w_sum_one_range9418w(0) <= sum_one(33);
	wire_tbl3_taylor_prod_w_sum_one_range9428w(0) <= sum_one(34);
	wire_tbl3_taylor_prod_w_sum_one_range9438w(0) <= sum_one(35);
	wire_tbl3_taylor_prod_w_sum_one_range9448w(0) <= sum_one(36);
	wire_tbl3_taylor_prod_w_sum_one_range9458w(0) <= sum_one(37);
	wire_tbl3_taylor_prod_w_sum_one_range9468w(0) <= sum_one(38);
	wire_tbl3_taylor_prod_w_sum_one_range9478w(0) <= sum_one(39);
	wire_tbl3_taylor_prod_w_sum_one_range9118w(0) <= sum_one(3);
	wire_tbl3_taylor_prod_w_sum_one_range9488w(0) <= sum_one(40);
	wire_tbl3_taylor_prod_w_sum_one_range9498w(0) <= sum_one(41);
	wire_tbl3_taylor_prod_w_sum_one_range9508w(0) <= sum_one(42);
	wire_tbl3_taylor_prod_w_sum_one_range9518w(0) <= sum_one(43);
	wire_tbl3_taylor_prod_w_sum_one_range9528w(0) <= sum_one(44);
	wire_tbl3_taylor_prod_w_sum_one_range9538w(0) <= sum_one(45);
	wire_tbl3_taylor_prod_w_sum_one_range9548w(0) <= sum_one(46);
	wire_tbl3_taylor_prod_w_sum_one_range9558w(0) <= sum_one(47);
	wire_tbl3_taylor_prod_w_sum_one_range9568w(0) <= sum_one(48);
	wire_tbl3_taylor_prod_w_sum_one_range9578w(0) <= sum_one(49);
	wire_tbl3_taylor_prod_w_sum_one_range9128w(0) <= sum_one(4);
	wire_tbl3_taylor_prod_w_sum_one_range9588w(0) <= sum_one(50);
	wire_tbl3_taylor_prod_w_sum_one_range9598w(0) <= sum_one(51);
	wire_tbl3_taylor_prod_w_sum_one_range9608w(0) <= sum_one(52);
	wire_tbl3_taylor_prod_w_sum_one_range9618w(0) <= sum_one(53);
	wire_tbl3_taylor_prod_w_sum_one_range9628w(0) <= sum_one(54);
	wire_tbl3_taylor_prod_w_sum_one_range9638w(0) <= sum_one(55);
	wire_tbl3_taylor_prod_w_sum_one_range9648w(0) <= sum_one(56);
	wire_tbl3_taylor_prod_w_sum_one_range9658w(0) <= sum_one(57);
	wire_tbl3_taylor_prod_w_sum_one_range9668w(0) <= sum_one(58);
	wire_tbl3_taylor_prod_w_sum_one_range9678w(0) <= sum_one(59);
	wire_tbl3_taylor_prod_w_sum_one_range9138w(0) <= sum_one(5);
	wire_tbl3_taylor_prod_w_sum_one_range9688w(0) <= sum_one(60);
	wire_tbl3_taylor_prod_w_sum_one_range9698w(0) <= sum_one(61);
	wire_tbl3_taylor_prod_w_sum_one_range9708w(0) <= sum_one(62);
	wire_tbl3_taylor_prod_w_sum_one_range9718w(0) <= sum_one(63);
	wire_tbl3_taylor_prod_w_sum_one_range9728w(0) <= sum_one(64);
	wire_tbl3_taylor_prod_w_sum_one_range9738w(0) <= sum_one(65);
	wire_tbl3_taylor_prod_w_sum_one_range9748w(0) <= sum_one(66);
	wire_tbl3_taylor_prod_w_sum_one_range9758w(0) <= sum_one(67);
	wire_tbl3_taylor_prod_w_sum_one_range9768w(0) <= sum_one(68);
	wire_tbl3_taylor_prod_w_sum_one_range9778w(0) <= sum_one(69);
	wire_tbl3_taylor_prod_w_sum_one_range9148w(0) <= sum_one(6);
	wire_tbl3_taylor_prod_w_sum_one_range9788w(0) <= sum_one(70);
	wire_tbl3_taylor_prod_w_sum_one_range9798w(0) <= sum_one(71);
	wire_tbl3_taylor_prod_w_sum_one_range9808w(0) <= sum_one(72);
	wire_tbl3_taylor_prod_w_sum_one_range9818w(0) <= sum_one(73);
	wire_tbl3_taylor_prod_w_sum_one_range9828w(0) <= sum_one(74);
	wire_tbl3_taylor_prod_w_sum_one_range9838w(0) <= sum_one(75);
	wire_tbl3_taylor_prod_w_sum_one_range9848w(0) <= sum_one(76);
	wire_tbl3_taylor_prod_w_sum_one_range9858w(0) <= sum_one(77);
	wire_tbl3_taylor_prod_w_sum_one_range9868w(0) <= sum_one(78);
	wire_tbl3_taylor_prod_w_sum_one_range9878w(0) <= sum_one(79);
	wire_tbl3_taylor_prod_w_sum_one_range9158w(0) <= sum_one(7);
	wire_tbl3_taylor_prod_w_sum_one_range9888w(0) <= sum_one(80);
	wire_tbl3_taylor_prod_w_sum_one_range9898w(0) <= sum_one(81);
	wire_tbl3_taylor_prod_w_sum_one_range9908w(0) <= sum_one(82);
	wire_tbl3_taylor_prod_w_sum_one_range9918w(0) <= sum_one(83);
	wire_tbl3_taylor_prod_w_sum_one_range9928w(0) <= sum_one(84);
	wire_tbl3_taylor_prod_w_sum_one_range9938w(0) <= sum_one(85);
	wire_tbl3_taylor_prod_w_sum_one_range9948w(0) <= sum_one(86);
	wire_tbl3_taylor_prod_w_sum_one_range9958w(0) <= sum_one(87);
	wire_tbl3_taylor_prod_w_sum_one_range9968w(0) <= sum_one(88);
	wire_tbl3_taylor_prod_w_sum_one_range9978w(0) <= sum_one(89);
	wire_tbl3_taylor_prod_w_sum_one_range9168w(0) <= sum_one(8);
	wire_tbl3_taylor_prod_w_sum_one_range9178w(0) <= sum_one(9);
	wire_tbl3_taylor_prod_w_vector1_range9990w(0) <= vector1(0);
	wire_tbl3_taylor_prod_w_vector1_range10102w(0) <= vector1(10);
	wire_tbl3_taylor_prod_w_vector1_range10113w(0) <= vector1(11);
	wire_tbl3_taylor_prod_w_vector1_range10124w(0) <= vector1(12);
	wire_tbl3_taylor_prod_w_vector1_range10135w(0) <= vector1(13);
	wire_tbl3_taylor_prod_w_vector1_range10146w(0) <= vector1(14);
	wire_tbl3_taylor_prod_w_vector1_range10157w(0) <= vector1(15);
	wire_tbl3_taylor_prod_w_vector1_range10168w(0) <= vector1(16);
	wire_tbl3_taylor_prod_w_vector1_range10179w(0) <= vector1(17);
	wire_tbl3_taylor_prod_w_vector1_range10190w(0) <= vector1(18);
	wire_tbl3_taylor_prod_w_vector1_range10201w(0) <= vector1(19);
	wire_tbl3_taylor_prod_w_vector1_range10003w(0) <= vector1(1);
	wire_tbl3_taylor_prod_w_vector1_range10212w(0) <= vector1(20);
	wire_tbl3_taylor_prod_w_vector1_range10223w(0) <= vector1(21);
	wire_tbl3_taylor_prod_w_vector1_range10234w(0) <= vector1(22);
	wire_tbl3_taylor_prod_w_vector1_range10245w(0) <= vector1(23);
	wire_tbl3_taylor_prod_w_vector1_range10256w(0) <= vector1(24);
	wire_tbl3_taylor_prod_w_vector1_range10267w(0) <= vector1(25);
	wire_tbl3_taylor_prod_w_vector1_range10278w(0) <= vector1(26);
	wire_tbl3_taylor_prod_w_vector1_range10289w(0) <= vector1(27);
	wire_tbl3_taylor_prod_w_vector1_range10300w(0) <= vector1(28);
	wire_tbl3_taylor_prod_w_vector1_range10311w(0) <= vector1(29);
	wire_tbl3_taylor_prod_w_vector1_range10014w(0) <= vector1(2);
	wire_tbl3_taylor_prod_w_vector1_range10322w(0) <= vector1(30);
	wire_tbl3_taylor_prod_w_vector1_range10333w(0) <= vector1(31);
	wire_tbl3_taylor_prod_w_vector1_range10344w(0) <= vector1(32);
	wire_tbl3_taylor_prod_w_vector1_range10355w(0) <= vector1(33);
	wire_tbl3_taylor_prod_w_vector1_range10366w(0) <= vector1(34);
	wire_tbl3_taylor_prod_w_vector1_range10377w(0) <= vector1(35);
	wire_tbl3_taylor_prod_w_vector1_range10388w(0) <= vector1(36);
	wire_tbl3_taylor_prod_w_vector1_range10399w(0) <= vector1(37);
	wire_tbl3_taylor_prod_w_vector1_range10410w(0) <= vector1(38);
	wire_tbl3_taylor_prod_w_vector1_range10421w(0) <= vector1(39);
	wire_tbl3_taylor_prod_w_vector1_range10025w(0) <= vector1(3);
	wire_tbl3_taylor_prod_w_vector1_range10432w(0) <= vector1(40);
	wire_tbl3_taylor_prod_w_vector1_range10443w(0) <= vector1(41);
	wire_tbl3_taylor_prod_w_vector1_range10454w(0) <= vector1(42);
	wire_tbl3_taylor_prod_w_vector1_range10465w(0) <= vector1(43);
	wire_tbl3_taylor_prod_w_vector1_range10476w(0) <= vector1(44);
	wire_tbl3_taylor_prod_w_vector1_range10487w(0) <= vector1(45);
	wire_tbl3_taylor_prod_w_vector1_range10498w(0) <= vector1(46);
	wire_tbl3_taylor_prod_w_vector1_range10509w(0) <= vector1(47);
	wire_tbl3_taylor_prod_w_vector1_range10520w(0) <= vector1(48);
	wire_tbl3_taylor_prod_w_vector1_range10531w(0) <= vector1(49);
	wire_tbl3_taylor_prod_w_vector1_range10036w(0) <= vector1(4);
	wire_tbl3_taylor_prod_w_vector1_range10542w(0) <= vector1(50);
	wire_tbl3_taylor_prod_w_vector1_range10553w(0) <= vector1(51);
	wire_tbl3_taylor_prod_w_vector1_range10564w(0) <= vector1(52);
	wire_tbl3_taylor_prod_w_vector1_range10575w(0) <= vector1(53);
	wire_tbl3_taylor_prod_w_vector1_range10586w(0) <= vector1(54);
	wire_tbl3_taylor_prod_w_vector1_range10597w(0) <= vector1(55);
	wire_tbl3_taylor_prod_w_vector1_range10608w(0) <= vector1(56);
	wire_tbl3_taylor_prod_w_vector1_range10619w(0) <= vector1(57);
	wire_tbl3_taylor_prod_w_vector1_range10630w(0) <= vector1(58);
	wire_tbl3_taylor_prod_w_vector1_range10641w(0) <= vector1(59);
	wire_tbl3_taylor_prod_w_vector1_range10047w(0) <= vector1(5);
	wire_tbl3_taylor_prod_w_vector1_range10652w(0) <= vector1(60);
	wire_tbl3_taylor_prod_w_vector1_range10663w(0) <= vector1(61);
	wire_tbl3_taylor_prod_w_vector1_range10674w(0) <= vector1(62);
	wire_tbl3_taylor_prod_w_vector1_range10685w(0) <= vector1(63);
	wire_tbl3_taylor_prod_w_vector1_range10696w(0) <= vector1(64);
	wire_tbl3_taylor_prod_w_vector1_range10707w(0) <= vector1(65);
	wire_tbl3_taylor_prod_w_vector1_range10718w(0) <= vector1(66);
	wire_tbl3_taylor_prod_w_vector1_range10729w(0) <= vector1(67);
	wire_tbl3_taylor_prod_w_vector1_range10740w(0) <= vector1(68);
	wire_tbl3_taylor_prod_w_vector1_range10751w(0) <= vector1(69);
	wire_tbl3_taylor_prod_w_vector1_range10058w(0) <= vector1(6);
	wire_tbl3_taylor_prod_w_vector1_range10762w(0) <= vector1(70);
	wire_tbl3_taylor_prod_w_vector1_range10773w(0) <= vector1(71);
	wire_tbl3_taylor_prod_w_vector1_range10784w(0) <= vector1(72);
	wire_tbl3_taylor_prod_w_vector1_range10795w(0) <= vector1(73);
	wire_tbl3_taylor_prod_w_vector1_range10806w(0) <= vector1(74);
	wire_tbl3_taylor_prod_w_vector1_range10817w(0) <= vector1(75);
	wire_tbl3_taylor_prod_w_vector1_range10828w(0) <= vector1(76);
	wire_tbl3_taylor_prod_w_vector1_range10839w(0) <= vector1(77);
	wire_tbl3_taylor_prod_w_vector1_range10850w(0) <= vector1(78);
	wire_tbl3_taylor_prod_w_vector1_range10861w(0) <= vector1(79);
	wire_tbl3_taylor_prod_w_vector1_range10069w(0) <= vector1(7);
	wire_tbl3_taylor_prod_w_vector1_range10872w(0) <= vector1(80);
	wire_tbl3_taylor_prod_w_vector1_range10883w(0) <= vector1(81);
	wire_tbl3_taylor_prod_w_vector1_range10894w(0) <= vector1(82);
	wire_tbl3_taylor_prod_w_vector1_range10905w(0) <= vector1(83);
	wire_tbl3_taylor_prod_w_vector1_range10916w(0) <= vector1(84);
	wire_tbl3_taylor_prod_w_vector1_range10927w(0) <= vector1(85);
	wire_tbl3_taylor_prod_w_vector1_range10938w(0) <= vector1(86);
	wire_tbl3_taylor_prod_w_vector1_range10949w(0) <= vector1(87);
	wire_tbl3_taylor_prod_w_vector1_range10960w(0) <= vector1(88);
	wire_tbl3_taylor_prod_w_vector1_range10971w(0) <= vector1(89);
	wire_tbl3_taylor_prod_w_vector1_range10080w(0) <= vector1(8);
	wire_tbl3_taylor_prod_w_vector1_range10091w(0) <= vector1(9);
	wire_tbl3_taylor_prod_w_vector2_range9083w(0) <= vector2(0);
	wire_tbl3_taylor_prod_w_vector2_range9185w(0) <= vector2(10);
	wire_tbl3_taylor_prod_w_vector2_range9195w(0) <= vector2(11);
	wire_tbl3_taylor_prod_w_vector2_range9205w(0) <= vector2(12);
	wire_tbl3_taylor_prod_w_vector2_range9215w(0) <= vector2(13);
	wire_tbl3_taylor_prod_w_vector2_range9225w(0) <= vector2(14);
	wire_tbl3_taylor_prod_w_vector2_range9235w(0) <= vector2(15);
	wire_tbl3_taylor_prod_w_vector2_range9245w(0) <= vector2(16);
	wire_tbl3_taylor_prod_w_vector2_range9255w(0) <= vector2(17);
	wire_tbl3_taylor_prod_w_vector2_range9265w(0) <= vector2(18);
	wire_tbl3_taylor_prod_w_vector2_range9275w(0) <= vector2(19);
	wire_tbl3_taylor_prod_w_vector2_range9095w(0) <= vector2(1);
	wire_tbl3_taylor_prod_w_vector2_range9285w(0) <= vector2(20);
	wire_tbl3_taylor_prod_w_vector2_range9295w(0) <= vector2(21);
	wire_tbl3_taylor_prod_w_vector2_range9305w(0) <= vector2(22);
	wire_tbl3_taylor_prod_w_vector2_range9315w(0) <= vector2(23);
	wire_tbl3_taylor_prod_w_vector2_range9325w(0) <= vector2(24);
	wire_tbl3_taylor_prod_w_vector2_range9335w(0) <= vector2(25);
	wire_tbl3_taylor_prod_w_vector2_range9345w(0) <= vector2(26);
	wire_tbl3_taylor_prod_w_vector2_range9355w(0) <= vector2(27);
	wire_tbl3_taylor_prod_w_vector2_range9365w(0) <= vector2(28);
	wire_tbl3_taylor_prod_w_vector2_range9375w(0) <= vector2(29);
	wire_tbl3_taylor_prod_w_vector2_range9105w(0) <= vector2(2);
	wire_tbl3_taylor_prod_w_vector2_range9385w(0) <= vector2(30);
	wire_tbl3_taylor_prod_w_vector2_range9395w(0) <= vector2(31);
	wire_tbl3_taylor_prod_w_vector2_range9405w(0) <= vector2(32);
	wire_tbl3_taylor_prod_w_vector2_range9415w(0) <= vector2(33);
	wire_tbl3_taylor_prod_w_vector2_range9425w(0) <= vector2(34);
	wire_tbl3_taylor_prod_w_vector2_range9435w(0) <= vector2(35);
	wire_tbl3_taylor_prod_w_vector2_range9445w(0) <= vector2(36);
	wire_tbl3_taylor_prod_w_vector2_range9455w(0) <= vector2(37);
	wire_tbl3_taylor_prod_w_vector2_range9465w(0) <= vector2(38);
	wire_tbl3_taylor_prod_w_vector2_range9475w(0) <= vector2(39);
	wire_tbl3_taylor_prod_w_vector2_range9115w(0) <= vector2(3);
	wire_tbl3_taylor_prod_w_vector2_range9485w(0) <= vector2(40);
	wire_tbl3_taylor_prod_w_vector2_range9495w(0) <= vector2(41);
	wire_tbl3_taylor_prod_w_vector2_range9505w(0) <= vector2(42);
	wire_tbl3_taylor_prod_w_vector2_range9515w(0) <= vector2(43);
	wire_tbl3_taylor_prod_w_vector2_range9525w(0) <= vector2(44);
	wire_tbl3_taylor_prod_w_vector2_range9535w(0) <= vector2(45);
	wire_tbl3_taylor_prod_w_vector2_range9545w(0) <= vector2(46);
	wire_tbl3_taylor_prod_w_vector2_range9555w(0) <= vector2(47);
	wire_tbl3_taylor_prod_w_vector2_range9565w(0) <= vector2(48);
	wire_tbl3_taylor_prod_w_vector2_range9575w(0) <= vector2(49);
	wire_tbl3_taylor_prod_w_vector2_range9125w(0) <= vector2(4);
	wire_tbl3_taylor_prod_w_vector2_range9585w(0) <= vector2(50);
	wire_tbl3_taylor_prod_w_vector2_range9595w(0) <= vector2(51);
	wire_tbl3_taylor_prod_w_vector2_range9605w(0) <= vector2(52);
	wire_tbl3_taylor_prod_w_vector2_range9615w(0) <= vector2(53);
	wire_tbl3_taylor_prod_w_vector2_range9625w(0) <= vector2(54);
	wire_tbl3_taylor_prod_w_vector2_range9635w(0) <= vector2(55);
	wire_tbl3_taylor_prod_w_vector2_range9645w(0) <= vector2(56);
	wire_tbl3_taylor_prod_w_vector2_range9655w(0) <= vector2(57);
	wire_tbl3_taylor_prod_w_vector2_range9665w(0) <= vector2(58);
	wire_tbl3_taylor_prod_w_vector2_range9675w(0) <= vector2(59);
	wire_tbl3_taylor_prod_w_vector2_range9135w(0) <= vector2(5);
	wire_tbl3_taylor_prod_w_vector2_range9685w(0) <= vector2(60);
	wire_tbl3_taylor_prod_w_vector2_range9695w(0) <= vector2(61);
	wire_tbl3_taylor_prod_w_vector2_range9705w(0) <= vector2(62);
	wire_tbl3_taylor_prod_w_vector2_range9715w(0) <= vector2(63);
	wire_tbl3_taylor_prod_w_vector2_range9725w(0) <= vector2(64);
	wire_tbl3_taylor_prod_w_vector2_range9735w(0) <= vector2(65);
	wire_tbl3_taylor_prod_w_vector2_range9745w(0) <= vector2(66);
	wire_tbl3_taylor_prod_w_vector2_range9755w(0) <= vector2(67);
	wire_tbl3_taylor_prod_w_vector2_range9765w(0) <= vector2(68);
	wire_tbl3_taylor_prod_w_vector2_range9775w(0) <= vector2(69);
	wire_tbl3_taylor_prod_w_vector2_range9145w(0) <= vector2(6);
	wire_tbl3_taylor_prod_w_vector2_range9785w(0) <= vector2(70);
	wire_tbl3_taylor_prod_w_vector2_range9795w(0) <= vector2(71);
	wire_tbl3_taylor_prod_w_vector2_range9805w(0) <= vector2(72);
	wire_tbl3_taylor_prod_w_vector2_range9815w(0) <= vector2(73);
	wire_tbl3_taylor_prod_w_vector2_range9825w(0) <= vector2(74);
	wire_tbl3_taylor_prod_w_vector2_range9835w(0) <= vector2(75);
	wire_tbl3_taylor_prod_w_vector2_range9845w(0) <= vector2(76);
	wire_tbl3_taylor_prod_w_vector2_range9855w(0) <= vector2(77);
	wire_tbl3_taylor_prod_w_vector2_range9865w(0) <= vector2(78);
	wire_tbl3_taylor_prod_w_vector2_range9875w(0) <= vector2(79);
	wire_tbl3_taylor_prod_w_vector2_range9155w(0) <= vector2(7);
	wire_tbl3_taylor_prod_w_vector2_range9885w(0) <= vector2(80);
	wire_tbl3_taylor_prod_w_vector2_range9895w(0) <= vector2(81);
	wire_tbl3_taylor_prod_w_vector2_range9905w(0) <= vector2(82);
	wire_tbl3_taylor_prod_w_vector2_range9915w(0) <= vector2(83);
	wire_tbl3_taylor_prod_w_vector2_range9925w(0) <= vector2(84);
	wire_tbl3_taylor_prod_w_vector2_range9935w(0) <= vector2(85);
	wire_tbl3_taylor_prod_w_vector2_range9945w(0) <= vector2(86);
	wire_tbl3_taylor_prod_w_vector2_range9955w(0) <= vector2(87);
	wire_tbl3_taylor_prod_w_vector2_range9965w(0) <= vector2(88);
	wire_tbl3_taylor_prod_w_vector2_range9975w(0) <= vector2(89);
	wire_tbl3_taylor_prod_w_vector2_range9165w(0) <= vector2(8);
	wire_tbl3_taylor_prod_w_vector2_range9175w(0) <= vector2(9);
	sum :  ALTFP_EXa_altmult_opt_csa_lsf
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => car_two_wo,
		datab => sum_two_wo,
		result => wire_sum_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN car_two_adj_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN car_two_adj_reg0 <= car_two_adj;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg0 <= lowest_bits_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg1 <= lowest_bits_wi_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_bits_wi_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lowest_bits_wi_reg2 <= lowest_bits_wi_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lsb_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN lsb_prod_wi_reg0 <= lsb_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mid_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mid_prod_wi_reg0 <= mid_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN msb_prod_wi_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN msb_prod_wi_reg0 <= msb_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sum_two_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sum_two_reg0 <= sum_two;
			END IF;
		END IF;
	END PROCESS;
	wire_compress_a_dataa <= ( "0" & wire_a(60 DOWNTO 31));
	compress_a :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		cout => wire_compress_a_cout,
		dataa => wire_compress_a_dataa,
		datab => wire_a(30 DOWNTO 0),
		result => wire_compress_a_result
	  );
	wire_compress_b_dataa <= ( "000" & wire_b(58 DOWNTO 31));
	compress_b :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		cout => wire_compress_b_cout,
		dataa => wire_compress_b_dataa,
		datab => wire_b(30 DOWNTO 0),
		result => wire_compress_b_result
	  );
	lsb_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 31,
		LPM_WIDTHB => 31,
		LPM_WIDTHP => 62,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_a(30 DOWNTO 0),
		datab => wire_b(30 DOWNTO 0),
		result => wire_lsb_prod_result
	  );
	wire_mid_prod_dataa <= ( wire_compress_a_cout & wire_compress_a_result);
	wire_mid_prod_datab <= ( wire_compress_b_cout & wire_compress_b_result);
	mid_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 32,
		LPM_WIDTHB => 32,
		LPM_WIDTHP => 64,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_mid_prod_dataa,
		datab => wire_mid_prod_datab,
		result => wire_mid_prod_result
	  );
	wire_msb_prod_dataa <= ( "0" & wire_a(60 DOWNTO 31));
	msb_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 31,
		LPM_WIDTHB => 28,
		LPM_WIDTHP => 59,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => wire_msb_prod_dataa,
		datab => wire_b(58 DOWNTO 31),
		result => wire_msb_prod_result
	  );

 END RTL; --ALTFP_EXa_altmult_opt_95e

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 18 lpm_clshift 1 lpm_compare 3 lpm_mult 11 lpm_mux 3 mux21 224 reg 2890 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTFP_EXa_altfp_exp_iuc IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END ALTFP_EXa_altfp_exp_iuc;

 ARCHITECTURE RTL OF ALTFP_EXa_altfp_exp_iuc IS

	 SIGNAL  wire_man_prod_result	:	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_result	:	STD_LOGIC_VECTOR (121 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_datab	:	STD_LOGIC_VECTOR (58 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_result	:	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_23_pipes22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_23_pipes22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_0	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_1	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_10	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_11	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_12	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_13	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_14	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_15	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_16	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_17	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_18	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_2	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_3	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_4	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_5	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_6	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_7	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_8	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_9	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_dffe1	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_extra_ln2_dffe_11_w_lg_q259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 extra_ln2_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fraction_dffe1	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_24_pipes23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_24_pipes23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_24_pipes23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_overflow_dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_round_dffe15	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_pipe_dffe16	:	STD_LOGIC_VECTOR(62 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 round_up_dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_dffe_w_lg_q3430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sign_dffe_w_lg_q3416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 table_one_dffe12	:	STD_LOGIC_VECTOR(60 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 table_three_dffe12	:	STD_LOGIC_VECTOR(60 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 table_two_dffe12	:	STD_LOGIC_VECTOR(60 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_10_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_0	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_1	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_2	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_3	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_4	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_5	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_6	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xf_pl_dffe12	:	STD_LOGIC_VECTOR(59 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xf_pre_2_dffe10	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xf_pre_dffe9	:	STD_LOGIC_VECTOR(69 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xi_exp_value_dffe4	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xi_ln2_prod_dffe7	:	STD_LOGIC_VECTOR(80 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xi_prod_dffe3	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_minus_bias_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_minus_bias_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_minus_bias_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_w_lg_w_result_range3427w3428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_w_result_range3427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_lg_w_lg_w_result_range3417w3418w3419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_lg_w_result_range3417w3418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_lg_w_lg_w_lg_w_result_range3417w3418w3419w3420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_result_range3417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_invert_exp_value_dataa	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_invert_exp_value_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_invert_exp_value_w_result_range232w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_man_round_datab	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_man_round_result	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_one_minus_xf_dataa	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_one_minus_xf_result	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_x_fixed_minus_xiln2_datab	:	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  wire_x_fixed_minus_xiln2_result	:	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  wire_xf_minus_ln2_datab	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_xf_minus_ln2_result	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_xi_add_one_datab	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_xi_add_one_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_result	:	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  wire_distance_overflow_comp_agb	:	STD_LOGIC;
	 SIGNAL  wire_tbl1_compare_ageb	:	STD_LOGIC;
	 SIGNAL  wire_underflow_compare_agb	:	STD_LOGIC;
	 SIGNAL  wire_xi_ln2_prod_result	:	STD_LOGIC_VECTOR (80 DOWNTO 0);
	 SIGNAL  wire_xi_prod_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_table_one_data_2d	:	STD_LOGIC_2D(511 DOWNTO 0, 60 DOWNTO 0);
	 SIGNAL  wire_table_one_result	:	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  wire_table_three_data_2d	:	STD_LOGIC_2D(511 DOWNTO 0, 41 DOWNTO 0);
	 SIGNAL  wire_table_three_result	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_table_two_data_2d	:	STD_LOGIC_2D(511 DOWNTO 0, 50 DOWNTO 0);
	 SIGNAL  wire_table_two_result	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL	wire_cin_to_bias_dataout	:	STD_LOGIC;
	 SIGNAL	wire_exp_result_mux_prea_dataout	:	STD_LOGIC_VECTOR(10 DOWNTO 0);
	 SIGNAL  wire_exp_result_mux_prea_w_lg_dataout3626w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL	wire_exp_value_b4_biasa_dataout	:	STD_LOGIC_VECTOR(10 DOWNTO 0);
	 SIGNAL	wire_exp_value_selecta_dataout	:	STD_LOGIC_VECTOR(6 DOWNTO 0);
	 SIGNAL	wire_exp_value_to_compare_muxa_dataout	:	STD_LOGIC_VECTOR(10 DOWNTO 0);
	 SIGNAL	wire_exp_value_to_ln2a_dataout	:	STD_LOGIC_VECTOR(10 DOWNTO 0);
	 SIGNAL	wire_extra_ln2_muxa_dataout	:	STD_LOGIC_VECTOR(59 DOWNTO 0);
	 SIGNAL	wire_man_result_muxa_dataout	:	STD_LOGIC_VECTOR(51 DOWNTO 0);
	 SIGNAL	wire_xf_muxa_dataout	:	STD_LOGIC_VECTOR(59 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_prod_shifted3390w	:	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_prod_wire3389w	:	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  wire_w_lg_underflow_w3623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range10w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range13w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range16w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range19w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range22w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range25w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range28w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range31w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range34w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range37w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_all_one_w_range62w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3677w3678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3632w3633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3637w3638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3642w3643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3647w3648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3652w3653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3657w3658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3662w3663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3667w3668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3672w3673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3474w3475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3477w3478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3480w3481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3483w3484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3486w3487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3489w3490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3492w3493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3495w3496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3498w3499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3501w3502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3447w3448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3504w3505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3507w3508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3510w3511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3513w3514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3516w3517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3519w3520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3522w3523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3525w3526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3528w3529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3531w3532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3450w3451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3534w3535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3537w3538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3540w3541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3543w3544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3546w3547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3549w3550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3552w3553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3555w3556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3558w3559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3561w3562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3453w3454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3564w3565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3567w3568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3570w3571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3573w3574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3576w3577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3579w3580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3582w3583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3585w3586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3588w3589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3591w3592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3456w3457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3594w3595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3597w3598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3459w3460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3462w3463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3465w3466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3468w3469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range3471w3472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_underflow_w3623w3624w3625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_shifter_underflow3622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_infinity_wo3425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_nan_wo3424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_zero_wo3426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_underflow_w3436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_data_not_zero_w_range218w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_wo_range3384w3388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_underflow_w3623w3624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w3620w3621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_overflow_w3605w3606w3607w3608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w3620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_overflow_w3605w3606w3607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_barrel_shifter_underflow3618w3619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_overflow_w3611w3612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_overflow_w3605w3606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_shifter_underflow3618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_distance_overflow3429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_distance_overflow3438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_overflow_w3611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_overflow_w3605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range117w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range120w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range144w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range147w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range69w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range153w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range156w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range159w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range162w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range165w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range174w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range177w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range180w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range72w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range183w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range186w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range189w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range195w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range198w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range204w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range75w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range213w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range10w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range13w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range16w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range19w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range22w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range25w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range28w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range78w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range31w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range34w35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range37w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range81w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range84w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range87w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3677w3679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3632w3635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3637w3640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3642w3645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3647w3650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3652w3655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3657w3660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3662w3665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3667w3670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range3672w3675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range3406w3407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range3403w3404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range3400w3401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range3397w3398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  addr_val_more_than_one :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  barrel_shifter_data :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  barrel_shifter_distance :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  barrel_shifter_underflow :	STD_LOGIC;
	 SIGNAL  barrel_shifter_underflow_wi :	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  distance_overflow :	STD_LOGIC;
	 SIGNAL  distance_overflow_val_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  distance_overflow_wi :	STD_LOGIC;
	 SIGNAL  exp_bias :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_bias_all_ones_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_data_all_one_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_data_not_zero_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_invert :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_one :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_out_all_one_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_out_not_zero_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_result_out :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_result_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_value :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  exp_value_wi :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  exp_value_wo :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  exp_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  extra_ln2 :	STD_LOGIC;
	 SIGNAL  fraction :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  fraction_wi :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  fraction_wo :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  gnd_w :	STD_LOGIC;
	 SIGNAL  guard_bit :	STD_LOGIC;
	 SIGNAL  input_is_infinity_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinity_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_wo :	STD_LOGIC;
	 SIGNAL  input_is_zero_wi :	STD_LOGIC;
	 SIGNAL  input_is_zero_wo :	STD_LOGIC;
	 SIGNAL  ln2_w :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  man_data_not_zero_w :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  man_overflow :	STD_LOGIC;
	 SIGNAL  man_overflow_wi :	STD_LOGIC;
	 SIGNAL  man_overflow_wo :	STD_LOGIC;
	 SIGNAL  man_prod_result :	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  man_prod_shifted :	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  man_prod_wi :	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  man_prod_wire :	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  man_prod_wo :	STD_LOGIC_VECTOR (119 DOWNTO 0);
	 SIGNAL  man_result_all_ones :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  man_result_w :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  man_round_wi :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  man_round_wo :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  nan_w :	STD_LOGIC;
	 SIGNAL  negative_infinity :	STD_LOGIC;
	 SIGNAL  one_over_ln2_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  overflow_w :	STD_LOGIC;
	 SIGNAL  positive_infinity :	STD_LOGIC;
	 SIGNAL  result_pipe_wi :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  result_pipe_wo :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  result_underflow_w :	STD_LOGIC;
	 SIGNAL  round_bit :	STD_LOGIC;
	 SIGNAL  round_up :	STD_LOGIC;
	 SIGNAL  round_up_wi :	STD_LOGIC;
	 SIGNAL  round_up_wo :	STD_LOGIC;
	 SIGNAL  shifted_value :	STD_LOGIC;
	 SIGNAL  sign_w :	STD_LOGIC;
	 SIGNAL  sticky_bits :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  table_one_data :	STD_LOGIC_VECTOR (31231 DOWNTO 0);
	 SIGNAL  table_one_out :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  table_one_out_pl :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  table_three_data :	STD_LOGIC_VECTOR (21503 DOWNTO 0);
	 SIGNAL  table_three_out :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  table_three_out_pl :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  table_three_out_tmp :	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  table_two_data :	STD_LOGIC_VECTOR (26111 DOWNTO 0);
	 SIGNAL  table_two_out :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  table_two_out_pl :	STD_LOGIC_VECTOR (60 DOWNTO 0);
	 SIGNAL  table_two_out_tmp :	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  tbl1_compare_wi :	STD_LOGIC;
	 SIGNAL  tbl1_compare_wo :	STD_LOGIC;
	 SIGNAL  tbl1_tbl2_prod_wi :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  tbl1_tbl2_prod_wo :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  tbl3_taylor_prod_wi :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  tbl3_taylor_prod_wo :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  underflow_compare_val_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  underflow_w :	STD_LOGIC;
	 SIGNAL  x_fixed :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  xf :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  xf_pl :	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  xf_pre :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  xf_pre_2_wi :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  xf_pre_2_wo :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  xf_pre_wi :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  xf_pre_wo :	STD_LOGIC_VECTOR (69 DOWNTO 0);
	 SIGNAL  xi_exp_value :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  xi_exp_value_wi :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  xi_exp_value_wo :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  xi_ln2_prod_wi :	STD_LOGIC_VECTOR (80 DOWNTO 0);
	 SIGNAL  xi_ln2_prod_wo :	STD_LOGIC_VECTOR (80 DOWNTO 0);
	 SIGNAL  xi_prod_wi :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  xi_prod_wo :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_data_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range3674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range3676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range3672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_value_wo_range234w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_exp_value_wo_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_value_wo_range231w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range3406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range3403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range3400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range3397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_wo_range3384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range3473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range3471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range3395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range3399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range3402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range3405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_xf_pre_2_wo_range285w	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 SIGNAL  wire_w_xf_pre_wo_range279w	:	STD_LOGIC_VECTOR (59 DOWNTO 0);
	 COMPONENT  ALTFP_EXa_altmult_opt_v4e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		dataa	:	IN  STD_LOGIC_VECTOR(59 DOWNTO 0);
		datab	:	IN  STD_LOGIC_VECTOR(59 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(119 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ALTFP_EXa_altmult_opt_45e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		dataa	:	IN  STD_LOGIC_VECTOR(60 DOWNTO 0);
		datab	:	IN  STD_LOGIC_VECTOR(60 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(121 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ALTFP_EXa_altmult_opt_95e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		dataa	:	IN  STD_LOGIC_VECTOR(60 DOWNTO 0);
		datab	:	IN  STD_LOGIC_VECTOR(58 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(119 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 119 GENERATE 
		wire_w_lg_man_prod_shifted3390w(i) <= man_prod_shifted(i) AND wire_w_man_prod_wo_range3384w(0);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 119 GENERATE 
		wire_w_lg_man_prod_wire3389w(i) <= man_prod_wire(i) AND wire_w_lg_w_man_prod_wo_range3384w3388w(0);
	END GENERATE loop1;
	wire_w_lg_underflow_w3623w(0) <= underflow_w AND wire_w_lg_barrel_shifter_underflow3622w(0);
	wire_w_lg_w_data_range10w43w(0) <= wire_w_data_range10w(0) AND wire_w_exp_data_all_one_w_range41w(0);
	wire_w_lg_w_data_range13w45w(0) <= wire_w_data_range13w(0) AND wire_w_exp_data_all_one_w_range44w(0);
	wire_w_lg_w_data_range16w47w(0) <= wire_w_data_range16w(0) AND wire_w_exp_data_all_one_w_range46w(0);
	wire_w_lg_w_data_range19w49w(0) <= wire_w_data_range19w(0) AND wire_w_exp_data_all_one_w_range48w(0);
	wire_w_lg_w_data_range22w51w(0) <= wire_w_data_range22w(0) AND wire_w_exp_data_all_one_w_range50w(0);
	wire_w_lg_w_data_range25w53w(0) <= wire_w_data_range25w(0) AND wire_w_exp_data_all_one_w_range52w(0);
	wire_w_lg_w_data_range28w55w(0) <= wire_w_data_range28w(0) AND wire_w_exp_data_all_one_w_range54w(0);
	wire_w_lg_w_data_range31w57w(0) <= wire_w_data_range31w(0) AND wire_w_exp_data_all_one_w_range56w(0);
	wire_w_lg_w_data_range34w59w(0) <= wire_w_data_range34w(0) AND wire_w_exp_data_all_one_w_range58w(0);
	wire_w_lg_w_data_range37w61w(0) <= wire_w_data_range37w(0) AND wire_w_exp_data_all_one_w_range60w(0);
	wire_w_lg_w_exp_data_all_one_w_range62w221w(0) <= wire_w_exp_data_all_one_w_range62w(0) AND wire_w_lg_w_man_data_not_zero_w_range218w220w(0);
	wire_w_lg_w_exp_result_w_range3677w3678w(0) <= wire_w_exp_result_w_range3677w(0) AND wire_w_exp_out_all_one_w_range3674w(0);
	wire_w_lg_w_exp_result_w_range3632w3633w(0) <= wire_w_exp_result_w_range3632w(0) AND wire_w_exp_out_all_one_w_range3628w(0);
	wire_w_lg_w_exp_result_w_range3637w3638w(0) <= wire_w_exp_result_w_range3637w(0) AND wire_w_exp_out_all_one_w_range3634w(0);
	wire_w_lg_w_exp_result_w_range3642w3643w(0) <= wire_w_exp_result_w_range3642w(0) AND wire_w_exp_out_all_one_w_range3639w(0);
	wire_w_lg_w_exp_result_w_range3647w3648w(0) <= wire_w_exp_result_w_range3647w(0) AND wire_w_exp_out_all_one_w_range3644w(0);
	wire_w_lg_w_exp_result_w_range3652w3653w(0) <= wire_w_exp_result_w_range3652w(0) AND wire_w_exp_out_all_one_w_range3649w(0);
	wire_w_lg_w_exp_result_w_range3657w3658w(0) <= wire_w_exp_result_w_range3657w(0) AND wire_w_exp_out_all_one_w_range3654w(0);
	wire_w_lg_w_exp_result_w_range3662w3663w(0) <= wire_w_exp_result_w_range3662w(0) AND wire_w_exp_out_all_one_w_range3659w(0);
	wire_w_lg_w_exp_result_w_range3667w3668w(0) <= wire_w_exp_result_w_range3667w(0) AND wire_w_exp_out_all_one_w_range3664w(0);
	wire_w_lg_w_exp_result_w_range3672w3673w(0) <= wire_w_exp_result_w_range3672w(0) AND wire_w_exp_out_all_one_w_range3669w(0);
	wire_w_lg_w_man_round_wi_range3474w3475w(0) <= wire_w_man_round_wi_range3474w(0) AND wire_w_man_result_all_ones_range3473w(0);
	wire_w_lg_w_man_round_wi_range3477w3478w(0) <= wire_w_man_round_wi_range3477w(0) AND wire_w_man_result_all_ones_range3476w(0);
	wire_w_lg_w_man_round_wi_range3480w3481w(0) <= wire_w_man_round_wi_range3480w(0) AND wire_w_man_result_all_ones_range3479w(0);
	wire_w_lg_w_man_round_wi_range3483w3484w(0) <= wire_w_man_round_wi_range3483w(0) AND wire_w_man_result_all_ones_range3482w(0);
	wire_w_lg_w_man_round_wi_range3486w3487w(0) <= wire_w_man_round_wi_range3486w(0) AND wire_w_man_result_all_ones_range3485w(0);
	wire_w_lg_w_man_round_wi_range3489w3490w(0) <= wire_w_man_round_wi_range3489w(0) AND wire_w_man_result_all_ones_range3488w(0);
	wire_w_lg_w_man_round_wi_range3492w3493w(0) <= wire_w_man_round_wi_range3492w(0) AND wire_w_man_result_all_ones_range3491w(0);
	wire_w_lg_w_man_round_wi_range3495w3496w(0) <= wire_w_man_round_wi_range3495w(0) AND wire_w_man_result_all_ones_range3494w(0);
	wire_w_lg_w_man_round_wi_range3498w3499w(0) <= wire_w_man_round_wi_range3498w(0) AND wire_w_man_result_all_ones_range3497w(0);
	wire_w_lg_w_man_round_wi_range3501w3502w(0) <= wire_w_man_round_wi_range3501w(0) AND wire_w_man_result_all_ones_range3500w(0);
	wire_w_lg_w_man_round_wi_range3447w3448w(0) <= wire_w_man_round_wi_range3447w(0) AND wire_w_man_result_all_ones_range3445w(0);
	wire_w_lg_w_man_round_wi_range3504w3505w(0) <= wire_w_man_round_wi_range3504w(0) AND wire_w_man_result_all_ones_range3503w(0);
	wire_w_lg_w_man_round_wi_range3507w3508w(0) <= wire_w_man_round_wi_range3507w(0) AND wire_w_man_result_all_ones_range3506w(0);
	wire_w_lg_w_man_round_wi_range3510w3511w(0) <= wire_w_man_round_wi_range3510w(0) AND wire_w_man_result_all_ones_range3509w(0);
	wire_w_lg_w_man_round_wi_range3513w3514w(0) <= wire_w_man_round_wi_range3513w(0) AND wire_w_man_result_all_ones_range3512w(0);
	wire_w_lg_w_man_round_wi_range3516w3517w(0) <= wire_w_man_round_wi_range3516w(0) AND wire_w_man_result_all_ones_range3515w(0);
	wire_w_lg_w_man_round_wi_range3519w3520w(0) <= wire_w_man_round_wi_range3519w(0) AND wire_w_man_result_all_ones_range3518w(0);
	wire_w_lg_w_man_round_wi_range3522w3523w(0) <= wire_w_man_round_wi_range3522w(0) AND wire_w_man_result_all_ones_range3521w(0);
	wire_w_lg_w_man_round_wi_range3525w3526w(0) <= wire_w_man_round_wi_range3525w(0) AND wire_w_man_result_all_ones_range3524w(0);
	wire_w_lg_w_man_round_wi_range3528w3529w(0) <= wire_w_man_round_wi_range3528w(0) AND wire_w_man_result_all_ones_range3527w(0);
	wire_w_lg_w_man_round_wi_range3531w3532w(0) <= wire_w_man_round_wi_range3531w(0) AND wire_w_man_result_all_ones_range3530w(0);
	wire_w_lg_w_man_round_wi_range3450w3451w(0) <= wire_w_man_round_wi_range3450w(0) AND wire_w_man_result_all_ones_range3449w(0);
	wire_w_lg_w_man_round_wi_range3534w3535w(0) <= wire_w_man_round_wi_range3534w(0) AND wire_w_man_result_all_ones_range3533w(0);
	wire_w_lg_w_man_round_wi_range3537w3538w(0) <= wire_w_man_round_wi_range3537w(0) AND wire_w_man_result_all_ones_range3536w(0);
	wire_w_lg_w_man_round_wi_range3540w3541w(0) <= wire_w_man_round_wi_range3540w(0) AND wire_w_man_result_all_ones_range3539w(0);
	wire_w_lg_w_man_round_wi_range3543w3544w(0) <= wire_w_man_round_wi_range3543w(0) AND wire_w_man_result_all_ones_range3542w(0);
	wire_w_lg_w_man_round_wi_range3546w3547w(0) <= wire_w_man_round_wi_range3546w(0) AND wire_w_man_result_all_ones_range3545w(0);
	wire_w_lg_w_man_round_wi_range3549w3550w(0) <= wire_w_man_round_wi_range3549w(0) AND wire_w_man_result_all_ones_range3548w(0);
	wire_w_lg_w_man_round_wi_range3552w3553w(0) <= wire_w_man_round_wi_range3552w(0) AND wire_w_man_result_all_ones_range3551w(0);
	wire_w_lg_w_man_round_wi_range3555w3556w(0) <= wire_w_man_round_wi_range3555w(0) AND wire_w_man_result_all_ones_range3554w(0);
	wire_w_lg_w_man_round_wi_range3558w3559w(0) <= wire_w_man_round_wi_range3558w(0) AND wire_w_man_result_all_ones_range3557w(0);
	wire_w_lg_w_man_round_wi_range3561w3562w(0) <= wire_w_man_round_wi_range3561w(0) AND wire_w_man_result_all_ones_range3560w(0);
	wire_w_lg_w_man_round_wi_range3453w3454w(0) <= wire_w_man_round_wi_range3453w(0) AND wire_w_man_result_all_ones_range3452w(0);
	wire_w_lg_w_man_round_wi_range3564w3565w(0) <= wire_w_man_round_wi_range3564w(0) AND wire_w_man_result_all_ones_range3563w(0);
	wire_w_lg_w_man_round_wi_range3567w3568w(0) <= wire_w_man_round_wi_range3567w(0) AND wire_w_man_result_all_ones_range3566w(0);
	wire_w_lg_w_man_round_wi_range3570w3571w(0) <= wire_w_man_round_wi_range3570w(0) AND wire_w_man_result_all_ones_range3569w(0);
	wire_w_lg_w_man_round_wi_range3573w3574w(0) <= wire_w_man_round_wi_range3573w(0) AND wire_w_man_result_all_ones_range3572w(0);
	wire_w_lg_w_man_round_wi_range3576w3577w(0) <= wire_w_man_round_wi_range3576w(0) AND wire_w_man_result_all_ones_range3575w(0);
	wire_w_lg_w_man_round_wi_range3579w3580w(0) <= wire_w_man_round_wi_range3579w(0) AND wire_w_man_result_all_ones_range3578w(0);
	wire_w_lg_w_man_round_wi_range3582w3583w(0) <= wire_w_man_round_wi_range3582w(0) AND wire_w_man_result_all_ones_range3581w(0);
	wire_w_lg_w_man_round_wi_range3585w3586w(0) <= wire_w_man_round_wi_range3585w(0) AND wire_w_man_result_all_ones_range3584w(0);
	wire_w_lg_w_man_round_wi_range3588w3589w(0) <= wire_w_man_round_wi_range3588w(0) AND wire_w_man_result_all_ones_range3587w(0);
	wire_w_lg_w_man_round_wi_range3591w3592w(0) <= wire_w_man_round_wi_range3591w(0) AND wire_w_man_result_all_ones_range3590w(0);
	wire_w_lg_w_man_round_wi_range3456w3457w(0) <= wire_w_man_round_wi_range3456w(0) AND wire_w_man_result_all_ones_range3455w(0);
	wire_w_lg_w_man_round_wi_range3594w3595w(0) <= wire_w_man_round_wi_range3594w(0) AND wire_w_man_result_all_ones_range3593w(0);
	wire_w_lg_w_man_round_wi_range3597w3598w(0) <= wire_w_man_round_wi_range3597w(0) AND wire_w_man_result_all_ones_range3596w(0);
	wire_w_lg_w_man_round_wi_range3459w3460w(0) <= wire_w_man_round_wi_range3459w(0) AND wire_w_man_result_all_ones_range3458w(0);
	wire_w_lg_w_man_round_wi_range3462w3463w(0) <= wire_w_man_round_wi_range3462w(0) AND wire_w_man_result_all_ones_range3461w(0);
	wire_w_lg_w_man_round_wi_range3465w3466w(0) <= wire_w_man_round_wi_range3465w(0) AND wire_w_man_result_all_ones_range3464w(0);
	wire_w_lg_w_man_round_wi_range3468w3469w(0) <= wire_w_man_round_wi_range3468w(0) AND wire_w_man_result_all_ones_range3467w(0);
	wire_w_lg_w_man_round_wi_range3471w3472w(0) <= wire_w_man_round_wi_range3471w(0) AND wire_w_man_result_all_ones_range3470w(0);
	wire_w_lg_w_lg_w_lg_underflow_w3623w3624w3625w(0) <= NOT wire_w_lg_w_lg_underflow_w3623w3624w(0);
	wire_w_lg_barrel_shifter_underflow3622w(0) <= NOT barrel_shifter_underflow;
	wire_w_lg_input_is_infinity_wo3425w(0) <= NOT input_is_infinity_wo;
	wire_w_lg_input_is_nan_wo3424w(0) <= NOT input_is_nan_wo;
	wire_w_lg_input_is_zero_wo3426w(0) <= NOT input_is_zero_wo;
	wire_w_lg_underflow_w3436w(0) <= NOT underflow_w;
	wire_w_lg_w_man_data_not_zero_w_range218w220w(0) <= NOT wire_w_man_data_not_zero_w_range218w(0);
	wire_w_lg_w_man_prod_wo_range3384w3388w(0) <= NOT wire_w_man_prod_wo_range3384w(0);
	wire_w_lg_w_lg_underflow_w3623w3624w(0) <= wire_w_lg_underflow_w3623w(0) OR negative_infinity;
	wire_w_lg_w3620w3621w(0) <= wire_w3620w(0) OR positive_infinity;
	wire_w_lg_w_lg_w_lg_w_lg_overflow_w3605w3606w3607w3608w(0) <= wire_w_lg_w_lg_w_lg_overflow_w3605w3606w3607w(0) OR input_is_infinity_wo;
	wire_w3620w(0) <= wire_w_lg_w_lg_barrel_shifter_underflow3618w3619w(0) OR nan_w;
	wire_w_lg_w_lg_w_lg_overflow_w3605w3606w3607w(0) <= wire_w_lg_w_lg_overflow_w3605w3606w(0) OR input_is_zero_wo;
	wire_w_lg_w_lg_barrel_shifter_underflow3618w3619w(0) <= wire_w_lg_barrel_shifter_underflow3618w(0) OR input_is_zero_wo;
	wire_w_lg_w_lg_overflow_w3611w3612w(0) <= wire_w_lg_overflow_w3611w(0) OR positive_infinity;
	wire_w_lg_w_lg_overflow_w3605w3606w(0) <= wire_w_lg_overflow_w3605w(0) OR nan_w;
	wire_w_lg_barrel_shifter_underflow3618w(0) <= barrel_shifter_underflow OR overflow_w;
	wire_w_lg_distance_overflow3429w(0) <= distance_overflow OR wire_exp_value_add_bias_w_lg_w_result_range3427w3428w(0);
	wire_w_lg_distance_overflow3438w(0) <= distance_overflow OR wire_exp_value_add_bias_w_result_range3427w(0);
	wire_w_lg_overflow_w3611w(0) <= overflow_w OR nan_w;
	wire_w_lg_overflow_w3605w(0) <= overflow_w OR underflow_w;
	wire_w_lg_w_data_range93w94w(0) <= wire_w_data_range93w(0) OR wire_w_man_data_not_zero_w_range92w(0);
	wire_w_lg_w_data_range96w97w(0) <= wire_w_data_range96w(0) OR wire_w_man_data_not_zero_w_range95w(0);
	wire_w_lg_w_data_range99w100w(0) <= wire_w_data_range99w(0) OR wire_w_man_data_not_zero_w_range98w(0);
	wire_w_lg_w_data_range102w103w(0) <= wire_w_data_range102w(0) OR wire_w_man_data_not_zero_w_range101w(0);
	wire_w_lg_w_data_range105w106w(0) <= wire_w_data_range105w(0) OR wire_w_man_data_not_zero_w_range104w(0);
	wire_w_lg_w_data_range108w109w(0) <= wire_w_data_range108w(0) OR wire_w_man_data_not_zero_w_range107w(0);
	wire_w_lg_w_data_range111w112w(0) <= wire_w_data_range111w(0) OR wire_w_man_data_not_zero_w_range110w(0);
	wire_w_lg_w_data_range114w115w(0) <= wire_w_data_range114w(0) OR wire_w_man_data_not_zero_w_range113w(0);
	wire_w_lg_w_data_range117w118w(0) <= wire_w_data_range117w(0) OR wire_w_man_data_not_zero_w_range116w(0);
	wire_w_lg_w_data_range120w121w(0) <= wire_w_data_range120w(0) OR wire_w_man_data_not_zero_w_range119w(0);
	wire_w_lg_w_data_range66w67w(0) <= wire_w_data_range66w(0) OR wire_w_man_data_not_zero_w_range64w(0);
	wire_w_lg_w_data_range123w124w(0) <= wire_w_data_range123w(0) OR wire_w_man_data_not_zero_w_range122w(0);
	wire_w_lg_w_data_range126w127w(0) <= wire_w_data_range126w(0) OR wire_w_man_data_not_zero_w_range125w(0);
	wire_w_lg_w_data_range129w130w(0) <= wire_w_data_range129w(0) OR wire_w_man_data_not_zero_w_range128w(0);
	wire_w_lg_w_data_range132w133w(0) <= wire_w_data_range132w(0) OR wire_w_man_data_not_zero_w_range131w(0);
	wire_w_lg_w_data_range135w136w(0) <= wire_w_data_range135w(0) OR wire_w_man_data_not_zero_w_range134w(0);
	wire_w_lg_w_data_range138w139w(0) <= wire_w_data_range138w(0) OR wire_w_man_data_not_zero_w_range137w(0);
	wire_w_lg_w_data_range141w142w(0) <= wire_w_data_range141w(0) OR wire_w_man_data_not_zero_w_range140w(0);
	wire_w_lg_w_data_range144w145w(0) <= wire_w_data_range144w(0) OR wire_w_man_data_not_zero_w_range143w(0);
	wire_w_lg_w_data_range147w148w(0) <= wire_w_data_range147w(0) OR wire_w_man_data_not_zero_w_range146w(0);
	wire_w_lg_w_data_range150w151w(0) <= wire_w_data_range150w(0) OR wire_w_man_data_not_zero_w_range149w(0);
	wire_w_lg_w_data_range69w70w(0) <= wire_w_data_range69w(0) OR wire_w_man_data_not_zero_w_range68w(0);
	wire_w_lg_w_data_range153w154w(0) <= wire_w_data_range153w(0) OR wire_w_man_data_not_zero_w_range152w(0);
	wire_w_lg_w_data_range156w157w(0) <= wire_w_data_range156w(0) OR wire_w_man_data_not_zero_w_range155w(0);
	wire_w_lg_w_data_range159w160w(0) <= wire_w_data_range159w(0) OR wire_w_man_data_not_zero_w_range158w(0);
	wire_w_lg_w_data_range162w163w(0) <= wire_w_data_range162w(0) OR wire_w_man_data_not_zero_w_range161w(0);
	wire_w_lg_w_data_range165w166w(0) <= wire_w_data_range165w(0) OR wire_w_man_data_not_zero_w_range164w(0);
	wire_w_lg_w_data_range168w169w(0) <= wire_w_data_range168w(0) OR wire_w_man_data_not_zero_w_range167w(0);
	wire_w_lg_w_data_range171w172w(0) <= wire_w_data_range171w(0) OR wire_w_man_data_not_zero_w_range170w(0);
	wire_w_lg_w_data_range174w175w(0) <= wire_w_data_range174w(0) OR wire_w_man_data_not_zero_w_range173w(0);
	wire_w_lg_w_data_range177w178w(0) <= wire_w_data_range177w(0) OR wire_w_man_data_not_zero_w_range176w(0);
	wire_w_lg_w_data_range180w181w(0) <= wire_w_data_range180w(0) OR wire_w_man_data_not_zero_w_range179w(0);
	wire_w_lg_w_data_range72w73w(0) <= wire_w_data_range72w(0) OR wire_w_man_data_not_zero_w_range71w(0);
	wire_w_lg_w_data_range183w184w(0) <= wire_w_data_range183w(0) OR wire_w_man_data_not_zero_w_range182w(0);
	wire_w_lg_w_data_range186w187w(0) <= wire_w_data_range186w(0) OR wire_w_man_data_not_zero_w_range185w(0);
	wire_w_lg_w_data_range189w190w(0) <= wire_w_data_range189w(0) OR wire_w_man_data_not_zero_w_range188w(0);
	wire_w_lg_w_data_range192w193w(0) <= wire_w_data_range192w(0) OR wire_w_man_data_not_zero_w_range191w(0);
	wire_w_lg_w_data_range195w196w(0) <= wire_w_data_range195w(0) OR wire_w_man_data_not_zero_w_range194w(0);
	wire_w_lg_w_data_range198w199w(0) <= wire_w_data_range198w(0) OR wire_w_man_data_not_zero_w_range197w(0);
	wire_w_lg_w_data_range201w202w(0) <= wire_w_data_range201w(0) OR wire_w_man_data_not_zero_w_range200w(0);
	wire_w_lg_w_data_range204w205w(0) <= wire_w_data_range204w(0) OR wire_w_man_data_not_zero_w_range203w(0);
	wire_w_lg_w_data_range207w208w(0) <= wire_w_data_range207w(0) OR wire_w_man_data_not_zero_w_range206w(0);
	wire_w_lg_w_data_range210w211w(0) <= wire_w_data_range210w(0) OR wire_w_man_data_not_zero_w_range209w(0);
	wire_w_lg_w_data_range75w76w(0) <= wire_w_data_range75w(0) OR wire_w_man_data_not_zero_w_range74w(0);
	wire_w_lg_w_data_range213w214w(0) <= wire_w_data_range213w(0) OR wire_w_man_data_not_zero_w_range212w(0);
	wire_w_lg_w_data_range216w217w(0) <= wire_w_data_range216w(0) OR wire_w_man_data_not_zero_w_range215w(0);
	wire_w_lg_w_data_range10w11w(0) <= wire_w_data_range10w(0) OR wire_w_exp_data_not_zero_w_range8w(0);
	wire_w_lg_w_data_range13w14w(0) <= wire_w_data_range13w(0) OR wire_w_exp_data_not_zero_w_range12w(0);
	wire_w_lg_w_data_range16w17w(0) <= wire_w_data_range16w(0) OR wire_w_exp_data_not_zero_w_range15w(0);
	wire_w_lg_w_data_range19w20w(0) <= wire_w_data_range19w(0) OR wire_w_exp_data_not_zero_w_range18w(0);
	wire_w_lg_w_data_range22w23w(0) <= wire_w_data_range22w(0) OR wire_w_exp_data_not_zero_w_range21w(0);
	wire_w_lg_w_data_range25w26w(0) <= wire_w_data_range25w(0) OR wire_w_exp_data_not_zero_w_range24w(0);
	wire_w_lg_w_data_range28w29w(0) <= wire_w_data_range28w(0) OR wire_w_exp_data_not_zero_w_range27w(0);
	wire_w_lg_w_data_range78w79w(0) <= wire_w_data_range78w(0) OR wire_w_man_data_not_zero_w_range77w(0);
	wire_w_lg_w_data_range31w32w(0) <= wire_w_data_range31w(0) OR wire_w_exp_data_not_zero_w_range30w(0);
	wire_w_lg_w_data_range34w35w(0) <= wire_w_data_range34w(0) OR wire_w_exp_data_not_zero_w_range33w(0);
	wire_w_lg_w_data_range37w38w(0) <= wire_w_data_range37w(0) OR wire_w_exp_data_not_zero_w_range36w(0);
	wire_w_lg_w_data_range81w82w(0) <= wire_w_data_range81w(0) OR wire_w_man_data_not_zero_w_range80w(0);
	wire_w_lg_w_data_range84w85w(0) <= wire_w_data_range84w(0) OR wire_w_man_data_not_zero_w_range83w(0);
	wire_w_lg_w_data_range87w88w(0) <= wire_w_data_range87w(0) OR wire_w_man_data_not_zero_w_range86w(0);
	wire_w_lg_w_data_range90w91w(0) <= wire_w_data_range90w(0) OR wire_w_man_data_not_zero_w_range89w(0);
	wire_w_lg_w_exp_result_w_range3677w3679w(0) <= wire_w_exp_result_w_range3677w(0) OR wire_w_exp_out_not_zero_w_range3676w(0);
	wire_w_lg_w_exp_result_w_range3632w3635w(0) <= wire_w_exp_result_w_range3632w(0) OR wire_w_exp_out_not_zero_w_range3630w(0);
	wire_w_lg_w_exp_result_w_range3637w3640w(0) <= wire_w_exp_result_w_range3637w(0) OR wire_w_exp_out_not_zero_w_range3636w(0);
	wire_w_lg_w_exp_result_w_range3642w3645w(0) <= wire_w_exp_result_w_range3642w(0) OR wire_w_exp_out_not_zero_w_range3641w(0);
	wire_w_lg_w_exp_result_w_range3647w3650w(0) <= wire_w_exp_result_w_range3647w(0) OR wire_w_exp_out_not_zero_w_range3646w(0);
	wire_w_lg_w_exp_result_w_range3652w3655w(0) <= wire_w_exp_result_w_range3652w(0) OR wire_w_exp_out_not_zero_w_range3651w(0);
	wire_w_lg_w_exp_result_w_range3657w3660w(0) <= wire_w_exp_result_w_range3657w(0) OR wire_w_exp_out_not_zero_w_range3656w(0);
	wire_w_lg_w_exp_result_w_range3662w3665w(0) <= wire_w_exp_result_w_range3662w(0) OR wire_w_exp_out_not_zero_w_range3661w(0);
	wire_w_lg_w_exp_result_w_range3667w3670w(0) <= wire_w_exp_result_w_range3667w(0) OR wire_w_exp_out_not_zero_w_range3666w(0);
	wire_w_lg_w_exp_result_w_range3672w3675w(0) <= wire_w_exp_result_w_range3672w(0) OR wire_w_exp_out_not_zero_w_range3671w(0);
	wire_w_lg_w_man_prod_result_range3406w3407w(0) <= wire_w_man_prod_result_range3406w(0) OR wire_w_sticky_bits_range3405w(0);
	wire_w_lg_w_man_prod_result_range3403w3404w(0) <= wire_w_man_prod_result_range3403w(0) OR wire_w_sticky_bits_range3402w(0);
	wire_w_lg_w_man_prod_result_range3400w3401w(0) <= wire_w_man_prod_result_range3400w(0) OR wire_w_sticky_bits_range3399w(0);
	wire_w_lg_w_man_prod_result_range3397w3398w(0) <= wire_w_man_prod_result_range3397w(0) OR wire_w_sticky_bits_range3395w(0);
	addr_val_more_than_one <= "101100011";
	barrel_shifter_data <= ( "00000000000" & "1" & fraction_wo & "000000");
	barrel_shifter_distance <= wire_exp_value_selecta_dataout;
	barrel_shifter_underflow <= barrel_shifter_underflow_dffe2_23_pipes22;
	barrel_shifter_underflow_wi <= (wire_underflow_compare_agb AND exp_value_wo(11));
	clk_en <= '1';
	distance_overflow <= distance_overflow_dffe2_23_pipes22;
	distance_overflow_val_w <= "00000001001";
	distance_overflow_wi <= (wire_distance_overflow_comp_agb AND (NOT exp_value_wo(11)));
	exp_bias <= "01111111111";
	exp_bias_all_ones_w <= (OTHERS => '1');
	exp_data_all_one_w <= ( wire_w_lg_w_data_range37w61w & wire_w_lg_w_data_range34w59w & wire_w_lg_w_data_range31w57w & wire_w_lg_w_data_range28w55w & wire_w_lg_w_data_range25w53w & wire_w_lg_w_data_range22w51w & wire_w_lg_w_data_range19w49w & wire_w_lg_w_data_range16w47w & wire_w_lg_w_data_range13w45w & wire_w_lg_w_data_range10w43w & data(52));
	exp_data_not_zero_w <= ( wire_w_lg_w_data_range37w38w & wire_w_lg_w_data_range34w35w & wire_w_lg_w_data_range31w32w & wire_w_lg_w_data_range28w29w & wire_w_lg_w_data_range25w26w & wire_w_lg_w_data_range22w23w & wire_w_lg_w_data_range19w20w & wire_w_lg_w_data_range16w17w & wire_w_lg_w_data_range13w14w & wire_w_lg_w_data_range10w11w & data(52));
	exp_invert <= (xi_exp_value XOR exp_bias_all_ones_w);
	exp_one <= ( wire_w_lg_w_lg_overflow_w3611w3612w & "1111111111");
	exp_out_all_one_w <= ( wire_w_lg_w_exp_result_w_range3677w3678w & wire_w_lg_w_exp_result_w_range3672w3673w & wire_w_lg_w_exp_result_w_range3667w3668w & wire_w_lg_w_exp_result_w_range3662w3663w & wire_w_lg_w_exp_result_w_range3657w3658w & wire_w_lg_w_exp_result_w_range3652w3653w & wire_w_lg_w_exp_result_w_range3647w3648w & wire_w_lg_w_exp_result_w_range3642w3643w & wire_w_lg_w_exp_result_w_range3637w3638w & wire_w_lg_w_exp_result_w_range3632w3633w & exp_result_w(0));
	exp_out_not_zero_w <= ( wire_w_lg_w_exp_result_w_range3677w3679w & wire_w_lg_w_exp_result_w_range3672w3675w & wire_w_lg_w_exp_result_w_range3667w3670w & wire_w_lg_w_exp_result_w_range3662w3665w & wire_w_lg_w_exp_result_w_range3657w3660w & wire_w_lg_w_exp_result_w_range3652w3655w & wire_w_lg_w_exp_result_w_range3647w3650w & wire_w_lg_w_exp_result_w_range3642w3645w & wire_w_lg_w_exp_result_w_range3637w3640w & wire_w_lg_w_exp_result_w_range3632w3635w & exp_result_w(0));
	exp_result_out <= wire_exp_result_mux_prea_w_lg_dataout3626w;
	exp_result_w <= wire_exp_value_man_over_result(10 DOWNTO 0);
	exp_value <= wire_exp_minus_bias_result;
	exp_value_wi <= exp_value;
	exp_value_wo <= exp_value_dffe1;
	exp_w <= data(62 DOWNTO 52);
	extra_ln2 <= ((NOT xf_pre(69)) AND sign_dffe10);
	fraction <= ( data(51 DOWNTO 0));
	fraction_wi <= fraction;
	fraction_wo <= fraction_dffe1;
	gnd_w <= '0';
	guard_bit <= man_prod_result(64);
	input_is_infinity_wi <= wire_w_lg_w_exp_data_all_one_w_range62w221w(0);
	input_is_infinity_wo <= input_is_infinity_24_pipes23;
	input_is_nan_wi <= (exp_data_all_one_w(10) AND man_data_not_zero_w(51));
	input_is_nan_wo <= input_is_nan_24_pipes23;
	input_is_zero_wi <= (NOT exp_data_not_zero_w(10));
	input_is_zero_wo <= input_is_zero_24_pipes23;
	ln2_w <= "1011000101110010000101111111011111010001110011110111100110101011110010";
	man_data_not_zero_w <= ( wire_w_lg_w_data_range216w217w & wire_w_lg_w_data_range213w214w & wire_w_lg_w_data_range210w211w & wire_w_lg_w_data_range207w208w & wire_w_lg_w_data_range204w205w & wire_w_lg_w_data_range201w202w & wire_w_lg_w_data_range198w199w & wire_w_lg_w_data_range195w196w & wire_w_lg_w_data_range192w193w & wire_w_lg_w_data_range189w190w & wire_w_lg_w_data_range186w187w & wire_w_lg_w_data_range183w184w & wire_w_lg_w_data_range180w181w & wire_w_lg_w_data_range177w178w & wire_w_lg_w_data_range174w175w & wire_w_lg_w_data_range171w172w & wire_w_lg_w_data_range168w169w & wire_w_lg_w_data_range165w166w & wire_w_lg_w_data_range162w163w & wire_w_lg_w_data_range159w160w & wire_w_lg_w_data_range156w157w & wire_w_lg_w_data_range153w154w & wire_w_lg_w_data_range150w151w & wire_w_lg_w_data_range147w148w & wire_w_lg_w_data_range144w145w & wire_w_lg_w_data_range141w142w & wire_w_lg_w_data_range138w139w & wire_w_lg_w_data_range135w136w & wire_w_lg_w_data_range132w133w & wire_w_lg_w_data_range129w130w & wire_w_lg_w_data_range126w127w & wire_w_lg_w_data_range123w124w & wire_w_lg_w_data_range120w121w & wire_w_lg_w_data_range117w118w & wire_w_lg_w_data_range114w115w & wire_w_lg_w_data_range111w112w & wire_w_lg_w_data_range108w109w & wire_w_lg_w_data_range105w106w & wire_w_lg_w_data_range102w103w & wire_w_lg_w_data_range99w100w & wire_w_lg_w_data_range96w97w & wire_w_lg_w_data_range93w94w & wire_w_lg_w_data_range90w91w & wire_w_lg_w_data_range87w88w & wire_w_lg_w_data_range84w85w & wire_w_lg_w_data_range81w82w & wire_w_lg_w_data_range78w79w & wire_w_lg_w_data_range75w76w & wire_w_lg_w_data_range72w73w & wire_w_lg_w_data_range69w70w & wire_w_lg_w_data_range66w67w & data(0));
	man_overflow <= (round_up AND man_result_all_ones(51));
	man_overflow_wi <= man_overflow;
	man_overflow_wo <= man_overflow_dffe15;
	man_prod_result <= (wire_w_lg_man_prod_shifted3390w OR wire_w_lg_man_prod_wire3389w);
	man_prod_shifted <= ( gnd_w & man_prod_wo(119 DOWNTO 1));
	man_prod_wi <= wire_man_prod_result;
	man_prod_wire <= man_prod_wo;
	man_prod_wo <= man_prod_wi;
	man_result_all_ones <= ( wire_w_lg_w_man_round_wi_range3597w3598w & wire_w_lg_w_man_round_wi_range3594w3595w & wire_w_lg_w_man_round_wi_range3591w3592w & wire_w_lg_w_man_round_wi_range3588w3589w & wire_w_lg_w_man_round_wi_range3585w3586w & wire_w_lg_w_man_round_wi_range3582w3583w & wire_w_lg_w_man_round_wi_range3579w3580w & wire_w_lg_w_man_round_wi_range3576w3577w & wire_w_lg_w_man_round_wi_range3573w3574w & wire_w_lg_w_man_round_wi_range3570w3571w & wire_w_lg_w_man_round_wi_range3567w3568w & wire_w_lg_w_man_round_wi_range3564w3565w & wire_w_lg_w_man_round_wi_range3561w3562w & wire_w_lg_w_man_round_wi_range3558w3559w & wire_w_lg_w_man_round_wi_range3555w3556w & wire_w_lg_w_man_round_wi_range3552w3553w & wire_w_lg_w_man_round_wi_range3549w3550w & wire_w_lg_w_man_round_wi_range3546w3547w & wire_w_lg_w_man_round_wi_range3543w3544w & wire_w_lg_w_man_round_wi_range3540w3541w & wire_w_lg_w_man_round_wi_range3537w3538w & wire_w_lg_w_man_round_wi_range3534w3535w & wire_w_lg_w_man_round_wi_range3531w3532w & wire_w_lg_w_man_round_wi_range3528w3529w & wire_w_lg_w_man_round_wi_range3525w3526w & wire_w_lg_w_man_round_wi_range3522w3523w & wire_w_lg_w_man_round_wi_range3519w3520w & wire_w_lg_w_man_round_wi_range3516w3517w & wire_w_lg_w_man_round_wi_range3513w3514w & wire_w_lg_w_man_round_wi_range3510w3511w & wire_w_lg_w_man_round_wi_range3507w3508w & wire_w_lg_w_man_round_wi_range3504w3505w & wire_w_lg_w_man_round_wi_range3501w3502w & wire_w_lg_w_man_round_wi_range3498w3499w & wire_w_lg_w_man_round_wi_range3495w3496w & wire_w_lg_w_man_round_wi_range3492w3493w & wire_w_lg_w_man_round_wi_range3489w3490w & wire_w_lg_w_man_round_wi_range3486w3487w & wire_w_lg_w_man_round_wi_range3483w3484w & wire_w_lg_w_man_round_wi_range3480w3481w & wire_w_lg_w_man_round_wi_range3477w3478w & wire_w_lg_w_man_round_wi_range3474w3475w & wire_w_lg_w_man_round_wi_range3471w3472w & wire_w_lg_w_man_round_wi_range3468w3469w & wire_w_lg_w_man_round_wi_range3465w3466w & wire_w_lg_w_man_round_wi_range3462w3463w & wire_w_lg_w_man_round_wi_range3459w3460w & wire_w_lg_w_man_round_wi_range3456w3457w
 & wire_w_lg_w_man_round_wi_range3453w3454w & wire_w_lg_w_man_round_wi_range3450w3451w & wire_w_lg_w_man_round_wi_range3447w3448w & man_round_wi(0));
	man_result_w <= wire_man_result_muxa_dataout;
	man_round_wi <= man_prod_result(115 DOWNTO 64);
	man_round_wo <= man_round_dffe15;
	nan_w <= input_is_nan_wo;
	negative_infinity <= (sign_dffe23 AND input_is_infinity_wo);
	one_over_ln2_w <= "101110001010";
	overflow_w <= (((wire_sign_dffe_w_lg_q3416w(0) AND ((wire_w_lg_distance_overflow3438w(0) OR exp_out_all_one_w(10)) OR wire_exp_value_man_over_result(11))) AND wire_w_lg_underflow_w3436w(0)) AND wire_w_lg_input_is_nan_wo3424w(0));
	positive_infinity <= (wire_sign_dffe_w_lg_q3416w(0) AND input_is_infinity_wo);
	result <= ( "0" & result_pipe_wo);
	result_pipe_wi <= ( exp_result_out & man_result_w);
	result_pipe_wo <= result_pipe_dffe16;
	result_underflow_w <= ((NOT exp_out_not_zero_w(10)) AND wire_exp_value_man_over_w_lg_w_lg_w_lg_w_result_range3417w3418w3419w3420w(0));
	round_bit <= man_prod_result(63);
	round_up <= (round_bit AND (guard_bit OR sticky_bits(4)));
	round_up_wi <= round_up;
	round_up_wo <= round_up_dffe15;
	shifted_value <= (tbl1_compare_wo OR man_prod_wo(117));
	sign_w <= data(63);
	sticky_bits <= ( wire_w_lg_w_man_prod_result_range3406w3407w & wire_w_lg_w_man_prod_result_range3403w3404w & wire_w_lg_w_man_prod_result_range3400w3401w & wire_w_lg_w_man_prod_result_range3397w3398w & man_prod_result(62));
	table_one_data <= ( "1010110110100001011011011110100111100001100100011101100101101" & "1010110101001010101100101110001101111100110010100110001010000" & "1010110011110100001000110010111111000101101000101101100100011" & "1010110010011101101111101011100100011000001011011101101111110" & "1010110001000111100001010110100111011011010011010100110010000" & "1010101111110001011101110010110010000000101011001110100010011" & "1010101110011011100100111110101110000100101111001110011011010" & "1010101101000101110110111001000101101110101011001001010110101" & "1010101011110000010011100000100011010000011001001111110101011" & "1010101010011010111010110011110001000110100000111000010000110" & "1010101001000101101100110001011001111000010101001001010111101" & "1010100111110000101001011000001000010111110011100100110101001" & "1010100110011011110000100110100111100001100010110010000011011" & "1010100101000111000010011011100010011100110001001001000111010" & "1010100011110010011110110101100100011011010011011101111000000" & "1010100010011110000101110011011000111001100011101011010001100" & "1010100001001001110111010011101011011110011111011110101111101" & "1010011111110101110011010101000111111011100111000011110110010" & "1010011110100001111001110110011010001100111011110000000010001" & "1010011101001110001010110110001110011000111110101110100101000" & "1010011011111010100110010011010000110000101111101100101100101" & "1010011010100111001100001100001101101111101011100101110010110" & "1010011001010011111100011111110001111011101011001111111001110" & "1010011000000000110111001100101010000101000010001000010001011" & "1010010110101101111100010001100011000110011101000000001000000" & "1010010101011011001011101101001010000101000000101001100100111" & "1010010100001000100101011110001100010000001000100100101101000" & "1010010010110110001001100011010111000001100101101100110011001" & "1010010001100011110111111011010111111101011101000101110001000" & "1010010000010001110000100100111100110010000110101001101011101" & "1010001110111111110011011110110011011000001011110110100001111"
 & "1010001101101110000000100111101001110010100110011100000100101" & "1010001100011100010111111110001110001110011111001001111010000" & "1010001011001010111001100001001111000011001100011101101010100" & "1010001001111001100101001111011010110010010001010001011000011" & "1010001000101000011011000111100000000111011011101010000001000" & "1010000111010111011011001000001101111000100011100110001000110" & "1010000110000110100101010000010011000101101001101100110000101" & "1010000100110101111001011110011110111000110101111100010110101" & "1010000011100101010111110001100000100110010110011001111111101" & "1010000010010101000000001000000111101100011110000000101011101" & "1010000001000100110010100001000011110011100011010000110100001" & "1001111111110100101110111011000100101101111110111111110100100" & "1001111110100100110101010100111010011000001011000111111100000" & "1001111101010101000101101101010100111000100001011000001010111" & "1001111100000101100000000011000100011111011010000100011000001" & "1001111010110110000100010100111001100111001010110101100010001" & "1001111001100110110010100001100100110100000101011010001001000" & "1001111000010111101010100111110110110100010110010110110010111" & "1001110111001000101100100110100000100000000011110110111010000" & "1001110101111001111000011100010010111001001100011101100101000" & "1001110100101011001110000111111111001011100101110110101000100" & "1001110011011100101101101000010110101100111011100111110011101" & "1001110010001110010110111100001010111100101110000010000100101" & "1001110001000000001010000010001101100100010000110011001001110" & "1001101111110010000110111001010000010110101001110111001001011" & "1001101110100100001101100000000101010000110000001010010101100" & "1001101101010110011101110101011110011001001010011011001000111" & "1001101100001000110111111000001110000000001101111100001101010" & "1001101010111011011011100111000110011111111101010110101011111" & "1001101001101110001001000000111010011100000111011100100111011" & "1001101000100001000000000100011100100010000101111011011111111" &
 "1001100111010100000000110000011111101000111100001110111111111" & "1001100110000111001011000011110110110001010110010011110011100" & "1001100100111010011110111101010101000101100111011010101001011" & "1001100011101101111100011011101101111001101000111011011100111" & "1001100010100001100011011101110100101010111001001000101001110" & "1001100001010101010100000010011101000000011010000010101001110" & "1001100000001001001110001000011010101010110000001011011011111" & "1001011110111101010001101110100001100100000001011010010100110" & "1001011101110001011110110011100101101111110011101111111000011" & "1001011100100101110101010110011011011011001100001001111110011" & "1001011011011010010101010101110110111100101101010111111110110" & "1001011010001110111110110000101100110100010110101111001000011" & "1001011001000011110001100101110001101011100010111111000000111" & "1001010111111000101101110011111010010101000111000110001110011" & "1001010110101101110011011001111011101101010001000111001010001" & "1001010101100011000010010110101010111001100110111100111100111" & "1001010100011000011010101000111101001001000101010000100100001" & "1001010011001101111100001111100111110011111110001110000001011" & "1001010010000011100111001001100000011011111000011001110010010" & "1001010000111001011011010101011100101011101101100110010010011" & "1001001111101111011000110010010010010111101001101001100101110" & "1001001110100101011111011110110111011101001001010011001101101" & "1001001101011011101111011010000010000010111001000010000101010" & "1001001100010010001000100010101000011000110011111010101001001" & "1001001011001000101010110111100000111000000010011101000110100" & "1001001001111111010110010111100010000010111001011011110100111" & "1001001000110110001011000001100010100100111000110001111000000" & "1001000111101101001000110100011001010010101010011001101011101" & "1001000110100100001111101110111101001010000001000011111000000" & "1001000101011011011111110000000101010001110111001110001111110" & "1001000100010010111000110110101000111010001101111010110110110" & "1001000011001010011011000001011111011100001011100111010010000"
 & "1001000010000010000110001111100000011001111011000100000001000" & "1001000000111001111010011111100011011110101010001011111111111" & "1000111111110001110111110000100000011110101000111100010010010" & "1000111110101001111110000001001111010111001000001011111000000" & "1000111101100010001101010000101000001110011000100011101010001" & "1000111100011010100101011101100011010011101001010110100001000" & "1000111011010011000110100110111000111111000111011001100100000" & "1000111010001011110000101011100001110001111011111100100001011" & "1000111001000100100011101010010110010110001011100010001111011" & "1000110111111101011111100010001111011110110100111001010110101" & "1000110110110110100100010010000110000111101111110101000100110" & "1000110101101111110001111000110011010101101100000110001000010" & "1000110100101001001000010101010000010110010000010011110101101" & "1000110011100010100111100110010110011111111000110101010100101" & "1000110010011100001111101010111111010001110110101010110110111" & "1000110001010110000000100010000100010100001110010111010111000" & "1000110000001111111010001010011111010111110110111010000000101" & "1000101111001001111100100011001010010110011000101000000001110" & "1000101110000100000111101010111111010010001100000110100011101" & "1000101100111110011011100000111000010110011001000100101101110" & "1000101011111000111000000011101111110110110101010101110000100" & "1000101010110011011101010010100000010000000011101011011001100" & "1000101001101110001011001100000100000111010010110000001111110" & "1000101000101001000001101111010110001010011100000010011000110" & "1000100111100100000000111011010001010000000010101110000111001" & "1000100110011111001000101110110000010111010010101000110000011" & "1000100101011010011001001000101110100111111111001011101100010" & "1000100100010101110010001000000111010010100010001111011100111" & "1000100011010001010011101011110101101111111011000110111111000" & "1000100010001100111101110010110101100001101101011011000010101" & "1000100001001000110000011100000010010010000000000101101101001" &
 "1000100000000100101011100110010111110011011100001110000011001" & "1000011111000000101111010000110010000001001100000011111010110" & "1000011101111100111011011010001100111110111001111011110111101" & "1000011100111001010000000001100100111000101111001011001101101" & "1000011011110101101101000101110110000011010011000100001101110" & "1000011010110010010010100101111100111011101001110010011010011" & "1000011001101111000000100000110110000111010011010111000100001" & "1000011000101011110110110101011110010100001010100101110000000" & "1000010111101000110101100010110010011000100100000001000100101" & "1000010110100101111100100111101111010011001100110111100000111" & "1000010101100011001100000011010010001011001010000000011010110" & "1000010100100000100011110100011000001111110110111001000110010" & "1000010011011110000011111001111110111001000100100010000100100" & "1000010010011011101100010011000011100110111000011100011100010" & "1000010001011001011100111110100100000001101011100111011001001" & "1000010000010111010101111011011101111010001001011101110100111" & "1000001111010101010111001000101111001001001110110100000111011" & "1000001110010011100000100101010101110000001000110101111111101" & "1000001101010001110010010000001111111000010100000100100101011" & "1000001100010000001100001000011011110011011011010100100010100" & "1000001011001110101110001100110111111011010110101100010011111" & "1000001010001101011000011100100010110010001010100010100100101" & "1000001001001100001010110110011011000010000110011100101110111" & "1000001000001011000101011001011111011101100100001101100110110" & "1000000111001010001000000100101110111111000110110100001100110" & "1000000110001001010010110111001000101001011001011010100111111" & "1000000101001000100101101111101011100111001110010101001000101" & "1000000100001000000000101101010111001011011110000001010011111" & "1000000011000111100011101111001010110001000110000101010101010" & "1000000010000111001110110100000101111011001000001111011010110" & "1000000001000111000001111011001000010100101001010101010111010" & "1000000000000110111101000011010001110000110000010100001110000"
 & "1111111110001110000000010111000100010101001010100000001010011" & "1111111100001110010110100101110011001010100000101000000011100" & "1111111010001110111100110000110000010111110001100100010011101" & "1111111000001111110010110101111100100011001000000111100000101" & "1111110110010000111000110011011000100010101001010011001111101" & "1111110100010010001110100111000101011100010010011000111011100" & "1111110010010011110100001111000100100101110110111010111010010" & "1111110000010101101001101001010111100100111110101101110011010" & "1111101110010111101110110100000000001111000011111010000100110" & "1111101100011010000011101101000000101001010000111101111001010" & "1111101010011100101000010010011011001000011110101111001100101" & "1111101000011111011100100010010010010001010010011110000001010" & "1111100110100010100000011010101000110111111011110111000100010" & "1111100100100101110011111001100010000000010011000110100010000" & "1111100010101001010110111101000000111101110110111011001001110" & "1111100000101101001001100011001001010011101010101001100001010" & "1111011110110001001011101001111110110100010100001111100111111" & "1111011100110101011101001111100101100001111010011000101001010" & "1111011010111001111110010010000001101110000010100000111111000" & "1111011000111110101110101111010111111001101110111010100010101" & "1111010111000011101110100101101100110101011100110001001110110" & "1111010101001000111101110011000101100001000010001111101110110" & "1111010011001110011100010101100111001011101100100100011111110" & "1111010001010100001010001011010111010011111110000110111110110" & "1111001111011010000111010010011011100111101100011101001000000" & "1111001101100000010011101000111010000011111110100001000100010" & "1111001011100110101111001100111000110101001010100111000110010" & "1111001001101101011001111100011110010110110100100011110110101" & "1111000111110100010011110101110001010011101011110010110000000" & "1111000101111011011100110110111000100101101001011100101001100" & "1111000100000010110100111101111011010101101110011110110000011" &
 "1111000010001010011100001001000000111100000001110001110001100" & "1111000000010010010010010110010000111111101110010001010000111" & "1110111110011010010111100011110011010111000001000011010001110" & "1110111100100010101011101111110000000111000111100000001011100" & "1110111010101011001110111000001111100100001101011010110000001" & "1110111000110100000000111011011010010001011011001000011111100" & "1110110110111101000001110111011001000000110011101010001011010" & "1110110101000110010001101010010100110011010010110100100111111" & "1110110011001111110000010010010110111000101011011001101110101" & "1110110001011001011101101101101000101111100101010001101100111" & "1110101111100011011001111010010100000101011011100100100010100" & "1110101101101101100100110110100010110110011010110011101111110" & "1110101011110111111110100000011111001101011111000100010001001" & "1110101010000010100110110110010011100100010010001000101010110" & "1110101000001101011101110110001010100011001001101011100001001" & "1110100110011000100011011110001111000001000101011010000010100" & "1110100100100011110111101100101100000011101101001110111101011" & "1110100010101111011010011111101100111111001111011101100110000" & "1110100000111011001011110101011101010110011110111101001010110" & "1110011111000111001011101100001000111010110001010100010110111" & "1110011101010011011010000001111011101011111101000101000100010" & "1110011011011111110110110101000001111000010111111000011010100" & "1110011001101100100010000011100111111100110100101010111101101" & "1110010111111001011011101011111010100100100001111001001011001" & "1110010110000110100011101100000110101001000111101100000100111" & "1110010100010011111010000010011001010010100110000110001010110" & "1110010010100001011110101100111111110111010011010000100010110" & "1110010000101111010001101010000111111011111001101000001111011" & "1110001110111101010010110111111111010011010110001011110100000" & "1110001101001011100010010100110011111110110110101001001000011" & "1110001011011001111111111110110100001101110111101011011001000" & "1110001001101000101011110100001110011110000011001001010111101"
 & "1110000111110111100101110011010001011011001110010011111000000" & "1110000110000110101101111010001011111111011000000100011100001" & "1110000100010110000100000111001101010010100111001100001110001" & "1110000010100101101000011000100100101011001000100011001000100" & "1110000000110101011010101100100001101101001101010111001100000" & "1101111111000101011011000001010100001011001001011100000100011" & "1101111101010101101001010101001100000101010001011010111010001" & "1101111011100110000101100110011001101001111001000010010011011" & "1101111001110110101111110011001101010101010001010110100001101" & "1101111000000111100111111001110111110001100111000001111110100" & "1101110110011000101101111000101001110111000000100101110101110" & "1101110100101010000001101101110100101011011100101010111101001" & "1101110010111011100011010111101001100010110000010010111010111" & "1101110001001101010010110100011001111110100101001001011000111" & "1101101111011111010000000010010111101110010111110101100111010" & "1101101101110001011010111111110100101111010110001100001010101" & "1101101100000011110011101011000011001100011101100000111010010" & "1101101010010110011010000010010101011110011000111001001010110" & "1101101000101001001110000011111110001011011111011110000110100" & "1101100110111100001111101110010000000111110010101111010100010" & "1101100101001111011110111111011110010100111100110101101011010" & "1101100011100010111011110101111100000010001110110110010100011" & "1101100001110110100110001111111100101100011111000101111010001" & "1101100000001010011110001011110011111110000111011100000100111" & "1101011110011110100011100111110101101111000011100111000101110" & "1101011100110010110110100010010110000100101111011111101101111" & "1101011011000111010110111001101001010010000101011101010100110" & "1101011001011100000100101100000011110111011100101010001010011" & "1101010111110000111111110111111010100010100111010111110111110" & "1101010110000110001000011011100010001110110001010100001101001" & "1101010100011011011110010101010000000100011101111101111100110" &
 "1101010010110001000001100011011001011001100110111010000011011" & "1101010001000110110010000100010011110001011010001000111110011" & "1101001111011100101111110110010100111100011000011100001111000" & "1101001101110010111010110111110010111000010011101100001010110" & "1101001100001001010011000111000011110000001101001101111001001" & "1101001010011111111000100010011101111100010100001001011110101" & "1101001000110110101011001000011000000010000011110000010101001" & "1101000111001101101010110111001000110100000001110011110001011" & "1101000101100100110111101101000111010001111100111011110101010" & "1101000011111100010001101000101010101000101010111110001111110" & "1101000010010011111000101000001010010010000111010101101001111" & "1101000000101011101100101001111101110101010001011001000000000" & "1100111111000011101101101100011101000110001010110011001010000" & "1100111101011011111011101110000000000101110101111010101101111" & "1100111011110100010110101100111111000010010100001010000010000" & "1100111010001100111110100111110010010110100100010111011010011" & "1100111000100101110011011100110010101010100001001101100011111" & "1100110110111110110101001010011000110010111111100100001100010" & "1100110101011000000011101110111101110001101100111000110110110" & "1100110011110001011111001000111010110101001101100111111110000" & "1100110010001011000111010110101001011000111011100110000010011" & "1100110000100100111100010110100011000101000100011001000101101" & "1100101110111110111110000111000001101110100111110010010011001" & "1100101101011001001100100110011111010111010110000111110100011" & "1100101011110011100111110011010110001101101110101110110011011" & "1100101010001110001111101100000000101100111110010101101000111" & "1100101000101001000100001110111001011100111101011110010111010" & "1100100111000100000101011010011011010010001110111001010011000" & "1100100101011111010011001101000001001101111101111111110110111" & "1100100011111010101101100101000110011101111101001111100100111" & "1100100010010110010100100001000110011100100100100101010100111" & "1100100000110010000111111111011100110000101111111000101101101"
 & "1100011111001110000111111110100101001101111101010111101101011" & "1100011101101010010100011100111011110100001100000010011011101" & "1100011100000110101101011000111100101111111010000111001010100" & "1100011010100011010010110001000100011010000011011110100010100" & "1100011001000000000100100011101111011000000000000111111011100" & "1100010111011101000010101111011010011011100010100110000010001" & "1100010101111010001101010010100010100010110110011011101010000" & "1100010100010111100100001011100100111000011110101000101011001" & "1100010010110101000111011000111110110011010100000111001101001" & "1100010001010010110110111001001101110110100100001000111101111" & "1100001111110000110010101010101111110001101110110100110100010" & "1100001110001110111010101100000010100000100101100100100000110" & "1100001100101101001110111011100100001011001001100010101000001" & "1100001011001011101111010111110011000101101010001000101011111" & "1100001001101010011011111111001101110000100011011101011110101" & "1100001000001001010100110000010010111000011100110011100100010" & "1100000110101000011001101001100001010110000111000111111110110" & "1100000101000111101010101001011000001110011011100001000110111" & "1100000011100111000111101110010110110010011001101101110001000" & "1100000010000110110000110110111100011111000110100100011110010" & "1100000000100110100110000001101000111101101010100010111001011" & "1011111111000110100111001100111100000011010000001101100000000" & "1011111101100110110100010111010101110001000010101111010111111" & "1011111100000111001101011111010110010100001100011010001111111" & "1011111010100111110010100011011110000101110101000110101101010" & "1011111001001000100011100010001101101011000000110100100100101" & "1011110111101001100000011010000101110100101110001011011111011" & "1011110110001010101001001001100111011111110100111011101100010" & "1011110100101011111101101111010011110101000100011110111100011" & "1011110011001101011110001001101100001001000010011001101100001" & "1011110001101111001010010111010001111100001000111100010111011" &
 "1011110000010001000010010110100110111010100101100100111010011" & "1011101110110011000110000110001100111100010111100000011101101" & "1011101101010101010101100100100110000101001110001101001101101" & "1011101011110111110000110000010100100100100111111100011111011" & "1011101010011010010111100111111010110101110000010100111111010" & "1011101000111101001010001001111011011111011110110101001100010" & "1011100111100000001000010100111001010100010101010101111110111" & "1011100110000011010010000111010111010010011110101101011011111" & "1011100100100110100111011111111000100011101101010001110010010" & "1011100011001010001000011101000000011101011001011100100101000" & "1011100001101101110100111101010010100000100000001110000000100" & "1011100000010001101100111111010010011001100001110000011011101" & "1011011110110101110000100001100100000000011111111100000100001" & "1011011101011001111111100010101011011000111100111010110110100" & "1011011011111110011010000001001100110001111001101100100001111" & "1011011010100010111111111011101100100101110100101010110110101" & "1011011001000111110001010000101111011010101000001110000001010" & "1011010111101100101101111110111010000001101001010001001111111" & "1011010110010001110110000100110001010111100101110111100100001" & "1011010100110111001001100000111010100100100011110000101111001" & "1011010011011100101000010001111010111011111110111110011010001" & "1011010010000010010010010110010111111100101000011001011001111" & "1011010000101000000111101100110111010000100100010111001101010" & "1011001111001110001000010011111110101101001001001111100111001" & "1011001101110100010100001010010100010010111110000010100100001" & "1011001100011010101011001110011110001101111000111110001011010" & "1011001011000001001101011111000010110100111110000100111001001" & "1011001001100111111010111010101000101010011101110011110111111" & "1011001000001110110011011111110110011011110011101001100000101" & "1011000110110101110111001101010011000001100100101100001001101" & "1011000101011101000110000001100101011111011110010000111110000" & "1011000100000100011111111011010101000100010100100011000010100"
 & "1011000010101100000100111001001001001010000001001010100011011" & "1011000001010011110100111001101001010101100001110100001110101" & "1010111111111011101111111011011101010110110110111000111001001" & "1010111110100011110101111101001101001001000010000101001110101" & "1010111101001100000110111101100000110010000101000001101100011" & "1010111011110100100010111011000000100010111111111010100111011" & "1010111010011101001001110100010100110111110000001000011101101" & "1010111001000101111011101000000110010111001110111000010001111" & "1010110111101110111000010100111101110011001111110100010010011" & "1010110110010111111111111001100100001000011111101100101010111" & "1010110101000001010010010100100010011110100011000000100001001" & "1010110011101010101111100100100010000111110100100110111100111" & "1010110010010100010111101000001100100001100100011000011001110" & "1010110000111110001010011110001011010011110101111000000100111" & "1010101111101000001000000101001000010001011110111101100100110" & "1010101110010010010000011011101101011000000110011110101100001" & "1010101100111100100011100000100100110000000010111001010111101" & "1010101011100111000001010010011000101100011000111101110110010" & "1010101010010001101001101111110011101010111010011000111100000" & "1010101000111100011100110111100000010100000100011110100000010" & "1010100111100111011010101000001001011010111110110100000101101" & "1010100110010010100011000000011001111101011001111011101101100" & "1010100100111101110101111110111101000011101101111110110101110" & "1010100011101001010011100010011110000000111001011001100001000" & "1010100010010100111011101001101000010010011111100101101001011" & "1010100001000000101110010011000111100000100111100110011110101" & "1010011111101100101011011101100111011101111010110100001101110" & "1010011110011000110011000111110100000111100011100111110011110" & "1010011101000101000101010000011001100101001100000110111010111" & "1010011011110001100001110110000100001000111100110000000010011" & "1010011010011110001000110111100000001111011011000110110000011" &
 "1010011001001010111010010011011010011111101000100000001110100" & "1010010111110111110110001000011111101011000000101111110001001" & "1010010110100100111100010101011100101101011000110011101000110" & "1010010101010010001100111000111110101100111101100001111101011" & "1010010011111111100111110001110010111010010010010101110101100" & "1010010010101101001100111110100110110000001111111100100101110" & "1010010001011010111100011110000111110100000011000011001100111" & "1010010000001000110110001111000011110101001011000011110111110" & "1010001110110110111010010000001000101101011000110011110001101" & "1010001101100101001000100000000100100000101101010000111101110" & "1010001100010011100000111101100101011101011000010000011011011" & "1010001011000010000011100111011001111011110111001100010011110" & "1010001001110000110000011100010000011110110011110010010011000" & "1010001000011111100111011010110111110011000010110010001010100" & "1010000111001110101000100001111110101111100010101100011101110" & "1010000101111101110011110000010100010101011010100001011001001" & "1010000100101101001001000100100111101111111000011111110011110" & "1010000011011100101000011101101000010100010000110100011001101" & "1010000010001100010001111010000101100001111100011001000001111" & "1010000000111100000101011000101111000010010111100100001101100" & "1001111111101100000010111000010100101001000000111000110001011" & "1001111110011100001010010111100110010011010111110101101001001" & "1001111101001100011011110101010100001000111011100101110101010" & "1001111011111100110111010000001110011011001001110000100001111" & "1001111010101101011100100111000101100101011101001001011001000" & "1001111001011110001011111000101010001101001100100000111101011" & "1001111000001111000101000011101101000001101001010101001111111" & "1001110111000000001000000110111110111011111110100010011111010" & "1001110101110001010101000001010000111111001111010100000000100" & "1001110100100010101011110001010100011000010101110101010010111" & "1001110011010100001100010101111010011110000010000011001011111" & "1001110010000101110110101101110100110000111000011101001110101"
 & "1001110000110111101010110111110100111011010000110111001100010" & "1001101111101001101000110010101100110001010101001010101110000" & "1001101110011011110000011101001110010001000000001001001001111" & "1001101101001110000001110110001011100001111100001101100000001" & "1001101100000000011100111100010110110101100010001110100011001" & "1001101010110011000001101110100010100110111000010001001000111" & "1001101001100101110000001011100001011010110000011010100101101" & "1001101000011000101000010010000101111111100111100011010001001" & "1001100111001011101010000001000011001101100100001001010101000" & "1001100101111110110101010111001100000110010101000011100100101" & "1001100100110010001010010011010011110101010000010100011111001" & "1001100011100101101000110100001101101111010001111101011010011" & "1001100010011001010000111000101101010010111010110001111000010" & "1001100001001101000010011111100110001000001111001011000101010" & "1001100000000000111101100111101100000000110101111011100000000" & "1001011110110101000010001111110010110111110111000010101011100" & "1001011101101001010000010110101110110001111010100001001001101" & "1001011100011101100111111011010011111101000111001100100000100" & "1001011011010010001000111100010110110001000001100011100111110" & "1001011010000110110011011000101011101110101010100011000000111" & "1001011000111011100111001111000111100000011110011001010111101" & "1001010111110000100100011110011110111010010011011100001100110" & "1001010110100101101011000101100110111001011000111100101010000" & "1001010101011010111011000011010100100100010101111100011110111" & "1001010100010000010100010110011101001011001000000011000111101" & "1001010011000101110110111101110110000111000010010010111101011" & "1001010001111011100010111000010100111010101011111110101110101" & "1001010000110001011000000100101111010001111111011111000010111" & "1001001111100111010110100001111011000010001001001000000101111" & "1001001110011101011110001110101110001001100101111111011100111" & "1001001101010011101111001001111110110000000010110010000101011" &
 "1001001100001010001001010010100011000110011010101010011100100" & "1001001011000000101100100111010001100110110110000110110000010" & "1001001001110111011001000111000000110100101001101111011001001" & "1001001000101110001110110000100111011100010101001101011110010" & "1001000111100101001101100010111100010011100010000001100000111" & "1001000110011100010101011100110110011001000010011010010010111" & "1001000101010011100110011101001100110100110000001011110101000" & "1001000100001011000000100010110110110111101011100110011111001" & "1001000011000010100011101100101011111011111010001110010001001" & "1001000001111010001111111001100011100100100101110010001100100" & "1001000000110010000101001000010101011101111011000011111000101" & "1000111111101010000011010111111001011101001000101111001101110" & "1000111110100010001010100111000111100000011110010010001011000" & "1000111101011010011010110100110111101111001010110100110100011" & "1000111100010010110100000000000010011001011100000001011001110" & "1000111011001011010110000111011111111000011100111100100111101" & "1000111010000100000001001010001000101110010100111101111111110" & "1000111000111100110101000110110101100110000110101000011011110" & "1000110111110101110001111100011111010011101110100010110111100" & "1000110110101110110111101001111110110100000010010001000110000" & "1000110101101000000110001110001101001100101111001100101101001" & "1000110100100001011101101000000011101100011001011110001100001" & "1000110011011010111101110110011011101010011010110110001010001" & "1000110010010100100110111000001110100111000001100110101101000" & "1000110001001110011000101100010110001011001111011100111010010" & "1000110000001000010011010001101100001000111000011010011111011" & "1000101111000010010110100111001010011010100001101111100100011" & "1000101101111100100010101011101011000011100000110100100101111" & "1000101100110110110111011110001000001111111010000100011000011" & "1000101011110001010100111101011100010100011111110110010100110" & "1000101010101011111011001000100001101110110001011000101100111" & "1000101001100110101001111110010011000100111001101011001000101"
 & "1000101000100001100001011101101011000101101110011001001100110" & "1000100111011100100001100101100100101000101110110101001001100" & "1000100110010111101010010100111010101110000010110010110001110" & "1000100101010010111011101010101000011110011001100010011011101" & "1000100100001110010101100101101001001011001000101100001000111" & "1000100011001001111000000100111000001110001011001010111000100" & "1000100010000101100011000111010001001010000000001000000000010" & "1000100001000001010110101011101111101001101001110110101111101" & "1000011111111101010010110001001111100000101100101111111010100" & "1000011110111001010111010110101100101011001110001101101101001" & "1000011101110101100100011011000011001101110011100111100111100" & "1000011100110001111001111101001111010101100001001110100010111" & "1000011011101110010111111100001101010111111001001000111101111" & "1000011010101010111110010110111001110010111010001111010010110" & "1000011001100111101101001100010001001100111111001000010101001" & "1000011000100100100100011011010000010100111101000101111000010" & "1000010111100001100100000010110100000010000011000001011110001" & "1000010110011110101100000001111001010011111000011001001110011" & "1000010101011011111100010111011101010010011100001100110110001" & "1000010100011001010101000010011101001110000011111010110000001" & "1000010011010110110110000001110110011111011010011101010100101" & "1000010010010100011111010100100110100111011111001000010010011" & "1000010001010010010000111001101011001111100100100110001111100" & "1000010000010000001010110000000010001001001111110110010011000" & "1000001111001110001100110110101001001110010111001001110110001" & "1000001110001100010111001100011110100001000001000010011101111" & "1000001101001010101001110000100000001011100011001111111110000" & "1000001100001001000100100001101100100000100001101110100010100" & "1000001011000111100111011111000001111010101101100101000010101" & "1000001010000110010010100111011110111101000100000011011011100" & "1000001001000101000101111010000010010010101101100001010010111" &
 "1000001000000100000001010101101010101110111100011100100010111" & "1000000111000011000100111001010111001101001100011000001100101" & "1000000110000010010000100100000110110001000000111011010100000" & "1000000101000001100100010100111000100110000100110000000011001" & "1000000100000001000000001010101100000000001000100010110110000" & "1000000011000000100100000100100000011011000010000001101110100" & "1000000010000000010000000001010101011010101010111011101111101" & "1000000001000000000100000000001010101011000000000000100010001" & "1000000000000000000000000000000000000000000000000000000000000");
	table_one_out <= wire_table_one_result;
	table_one_out_pl <= table_one_dffe12;
	table_three_data <= ( "111111111000000000011111111000000000101010" & "111111110000000000011111110000000010001010" & "111111101000000000011111101000000100101010" & "111111100000000000011111100000001000001010" & "111111011000000000011111011000001100101010" & "111111010000000000011111010000010010001010" & "111111001000000000011111001000011000101010" & "111111000000000000011111000000100000001010" & "111110111000000000011110111000101000101010" & "111110110000000000011110110000110010001010" & "111110101000000000011110101000111100101001" & "111110100000000000011110100001001000001001" & "111110011000000000011110011001010100101001" & "111110010000000000011110010001100010001001" & "111110001000000000011110001001110000101001" & "111110000000000000011110000010000000001001" & "111101111000000000011101111010010000101001" & "111101110000000000011101110010100010001001" & "111101101000000000011101101010110100101001" & "111101100000000000011101100011001000001001" & "111101011000000000011101011011011100101001" & "111101010000000000011101010011110010001001" & "111101001000000000011101001100001000101001" & "111101000000000000011101000100100000001001" & "111100111000000000011100111100111000101001" & "111100110000000000011100110101010010001001" & "111100101000000000011100101101101100101001" & "111100100000000000011100100110001000001001" & "111100011000000000011100011110100100101000" & "111100010000000000011100010111000010001000" & "111100001000000000011100001111100000101000" & "111100000000000000011100001000000000001000" & "111011111000000000011100000000100000101000" & "111011110000000000011011111001000010001000" & "111011101000000000011011110001100100101000" & "111011100000000000011011101010001000001000" & "111011011000000000011011100010101100101000" & "111011010000000000011011011011010010001000" & "111011001000000000011011010011111000101000" & "111011000000000000011011001100100000001000" & "111010111000000000011011000101001000101000" & "111010110000000000011010111101110010001000" & "111010101000000000011010110110011100101000" & "111010100000000000011010101111001000001000"
 & "111010011000000000011010100111110100101000" & "111010010000000000011010100000100010001000" & "111010001000000000011010011001010000100111" & "111010000000000000011010010010000000000111" & "111001111000000000011010001010110000100111" & "111001110000000000011010000011100010000111" & "111001101000000000011001111100010100100111" & "111001100000000000011001110101001000000111" & "111001011000000000011001101101111100100111" & "111001010000000000011001100110110010000111" & "111001001000000000011001011111101000100111" & "111001000000000000011001011000100000000111" & "111000111000000000011001010001011000100111" & "111000110000000000011001001010010010000111" & "111000101000000000011001000011001100100111" & "111000100000000000011000111100001000000111" & "111000011000000000011000110101000100100111" & "111000010000000000011000101110000010000111" & "111000001000000000011000100111000000100111" & "111000000000000000011000100000000000000111" & "110111111000000000011000011001000000100111" & "110111110000000000011000010010000010000111" & "110111101000000000011000001011000100100111" & "110111100000000000011000000100001000000110" & "110111011000000000010111111101001100100110" & "110111010000000000010111110110010010000110" & "110111001000000000010111101111011000100110" & "110111000000000000010111101000100000000110" & "110110111000000000010111100001101000100110" & "110110110000000000010111011010110010000110" & "110110101000000000010111010011111100100110" & "110110100000000000010111001101001000000110" & "110110011000000000010111000110010100100110" & "110110010000000000010110111111100010000110" & "110110001000000000010110111000110000100110" & "110110000000000000010110110010000000000110" & "110101111000000000010110101011010000100110" & "110101110000000000010110100100100010000110" & "110101101000000000010110011101110100100110" & "110101100000000000010110010111001000000110" & "110101011000000000010110010000011100100110" & "110101010000000000010110001001110010000110" & "110101001000000000010110000011001000100110" & "110101000000000000010101111100100000000110"
 & "110100111000000000010101110101111000100110" & "110100110000000000010101101111010010000101" & "110100101000000000010101101000101100100101" & "110100100000000000010101100010001000000101" & "110100011000000000010101011011100100100101" & "110100010000000000010101010101000010000101" & "110100001000000000010101001110100000100101" & "110100000000000000010101001000000000000101" & "110011111000000000010101000001100000100101" & "110011110000000000010100111011000010000101" & "110011101000000000010100110100100100100101" & "110011100000000000010100101110001000000101" & "110011011000000000010100100111101100100101" & "110011010000000000010100100001010010000101" & "110011001000000000010100011010111000100101" & "110011000000000000010100010100100000000101" & "110010111000000000010100001110001000100101" & "110010110000000000010100000111110010000101" & "110010101000000000010100000001011100100101" & "110010100000000000010011111011001000000101" & "110010011000000000010011110100110100100101" & "110010010000000000010011101110100010000101" & "110010001000000000010011101000010000100101" & "110010000000000000010011100010000000000101" & "110001111000000000010011011011110000100101" & "110001110000000000010011010101100010000101" & "110001101000000000010011001111010100100100" & "110001100000000000010011001001001000000100" & "110001011000000000010011000010111100100100" & "110001010000000000010010111100110010000100" & "110001001000000000010010110110101000100100" & "110001000000000000010010110000100000000100" & "110000111000000000010010101010011000100100" & "110000110000000000010010100100010010000100" & "110000101000000000010010011110001100100100" & "110000100000000000010010011000001000000100" & "110000011000000000010010010010000100100100" & "110000010000000000010010001100000010000100" & "110000001000000000010010000110000000100100" & "110000000000000000010010000000000000000100" & "101111111000000000010001111010000000100100" & "101111110000000000010001110100000010000100" & "101111101000000000010001101110000100100100" & "101111100000000000010001101000001000000100"
 & "101111011000000000010001100010001100100100" & "101111010000000000010001011100010010000100" & "101111001000000000010001010110011000100100" & "101111000000000000010001010000100000000100" & "101110111000000000010001001010101000100100" & "101110110000000000010001000100110010000100" & "101110101000000000010000111110111100100100" & "101110100000000000010000111001001000000100" & "101110011000000000010000110011010100100100" & "101110010000000000010000101101100010000100" & "101110001000000000010000100111110000100011" & "101110000000000000010000100010000000000011" & "101101111000000000010000011100010000100011" & "101101110000000000010000010110100010000011" & "101101101000000000010000010000110100100011" & "101101100000000000010000001011001000000011" & "101101011000000000010000000101011100100011" & "101101010000000000001111111111110010000011" & "101101001000000000001111111010001000100011" & "101101000000000000001111110100100000000011" & "101100111000000000001111101110111000100011" & "101100110000000000001111101001010010000011" & "101100101000000000001111100011101100100011" & "101100100000000000001111011110001000000011" & "101100011000000000001111011000100100100011" & "101100010000000000001111010011000010000011" & "101100001000000000001111001101100000100011" & "101100000000000000001111001000000000000011" & "101011111000000000001111000010100000100011" & "101011110000000000001110111101000010000011" & "101011101000000000001110110111100100100011" & "101011100000000000001110110010001000000011" & "101011011000000000001110101100101100100011" & "101011010000000000001110100111010010000011" & "101011001000000000001110100001111000100011" & "101011000000000000001110011100100000000011" & "101010111000000000001110010111001000100011" & "101010110000000000001110010001110010000011" & "101010101000000000001110001100011100100011" & "101010100000000000001110000111001000000011" & "101010011000000000001110000001110100100011" & "101010010000000000001101111100100010000011" & "101010001000000000001101110111010000100011" & "101010000000000000001101110010000000000011"
 & "101001111000000000001101101100110000100010" & "101001110000000000001101100111100010000010" & "101001101000000000001101100010010100100010" & "101001100000000000001101011101001000000010" & "101001011000000000001101010111111100100010" & "101001010000000000001101010010110010000010" & "101001001000000000001101001101101000100010" & "101001000000000000001101001000100000000010" & "101000111000000000001101000011011000100010" & "101000110000000000001100111110010010000010" & "101000101000000000001100111001001100100010" & "101000100000000000001100110100001000000010" & "101000011000000000001100101111000100100010" & "101000010000000000001100101010000010000010" & "101000001000000000001100100101000000100010" & "101000000000000000001100100000000000000010" & "100111111000000000001100011011000000100010" & "100111110000000000001100010110000010000010" & "100111101000000000001100010001000100100010" & "100111100000000000001100001100001000000010" & "100111011000000000001100000111001100100010" & "100111010000000000001100000010010010000010" & "100111001000000000001011111101011000100010" & "100111000000000000001011111000100000000010" & "100110111000000000001011110011101000100010" & "100110110000000000001011101110110010000010" & "100110101000000000001011101001111100100010" & "100110100000000000001011100101001000000010" & "100110011000000000001011100000010100100010" & "100110010000000000001011011011100010000010" & "100110001000000000001011010110110000100010" & "100110000000000000001011010010000000000010" & "100101111000000000001011001101010000100010" & "100101110000000000001011001000100010000010" & "100101101000000000001011000011110100100010" & "100101100000000000001010111111001000000010" & "100101011000000000001010111010011100100010" & "100101010000000000001010110101110010000010" & "100101001000000000001010110001001000100010" & "100101000000000000001010101100100000000010" & "100100111000000000001010100111111000100010" & "100100110000000000001010100011010010000010" & "100100101000000000001010011110101100100001" & "100100100000000000001010011010001000000001"
 & "100100011000000000001010010101100100100001" & "100100010000000000001010010001000010000001" & "100100001000000000001010001100100000100001" & "100100000000000000001010001000000000000001" & "100011111000000000001010000011100000100001" & "100011110000000000001001111111000010000001" & "100011101000000000001001111010100100100001" & "100011100000000000001001110110001000000001" & "100011011000000000001001110001101100100001" & "100011010000000000001001101101010010000001" & "100011001000000000001001101000111000100001" & "100011000000000000001001100100100000000001" & "100010111000000000001001100000001000100001" & "100010110000000000001001011011110010000001" & "100010101000000000001001010111011100100001" & "100010100000000000001001010011001000000001" & "100010011000000000001001001110110100100001" & "100010010000000000001001001010100010000001" & "100010001000000000001001000110010000100001" & "100010000000000000001001000010000000000001" & "100001111000000000001000111101110000100001" & "100001110000000000001000111001100010000001" & "100001101000000000001000110101010100100001" & "100001100000000000001000110001001000000001" & "100001011000000000001000101100111100100001" & "100001010000000000001000101000110010000001" & "100001001000000000001000100100101000100001" & "100001000000000000001000100000100000000001" & "100000111000000000001000011100011000100001" & "100000110000000000001000011000010010000001" & "100000101000000000001000010100001100100001" & "100000100000000000001000010000001000000001" & "100000011000000000001000001100000100100001" & "100000010000000000001000001000000010000001" & "100000001000000000001000000100000000100001" & "100000000000000000001000000000000000000001" & "011111111000000000000111111100000000100001" & "011111110000000000000111111000000010000001" & "011111101000000000000111110100000100100001" & "011111100000000000000111110000001000000001" & "011111011000000000000111101100001100100001" & "011111010000000000000111101000010010000001" & "011111001000000000000111100100011000100001" & "011111000000000000000111100000100000000001"
 & "011110111000000000000111011100101000100001" & "011110110000000000000111011000110010000001" & "011110101000000000000111010100111100100001" & "011110100000000000000111010001001000000001" & "011110011000000000000111001101010100100001" & "011110010000000000000111001001100010000001" & "011110001000000000000111000101110000100001" & "011110000000000000000111000010000000000001" & "011101111000000000000110111110010000100001" & "011101110000000000000110111010100010000001" & "011101101000000000000110110110110100100001" & "011101100000000000000110110011001000000001" & "011101011000000000000110101111011100100001" & "011101010000000000000110101011110010000001" & "011101001000000000000110101000001000100001" & "011101000000000000000110100100100000000000" & "011100111000000000000110100000111000100000" & "011100110000000000000110011101010010000000" & "011100101000000000000110011001101100100000" & "011100100000000000000110010110001000000000" & "011100011000000000000110010010100100100000" & "011100010000000000000110001111000010000000" & "011100001000000000000110001011100000100000" & "011100000000000000000110001000000000000000" & "011011111000000000000110000100100000100000" & "011011110000000000000110000001000010000000" & "011011101000000000000101111101100100100000" & "011011100000000000000101111010001000000000" & "011011011000000000000101110110101100100000" & "011011010000000000000101110011010010000000" & "011011001000000000000101101111111000100000" & "011011000000000000000101101100100000000000" & "011010111000000000000101101001001000100000" & "011010110000000000000101100101110010000000" & "011010101000000000000101100010011100100000" & "011010100000000000000101011111001000000000" & "011010011000000000000101011011110100100000" & "011010010000000000000101011000100010000000" & "011010001000000000000101010101010000100000" & "011010000000000000000101010010000000000000" & "011001111000000000000101001110110000100000" & "011001110000000000000101001011100010000000" & "011001101000000000000101001000010100100000" & "011001100000000000000101000101001000000000"
 & "011001011000000000000101000001111100100000" & "011001010000000000000100111110110010000000" & "011001001000000000000100111011101000100000" & "011001000000000000000100111000100000000000" & "011000111000000000000100110101011000100000" & "011000110000000000000100110010010010000000" & "011000101000000000000100101111001100100000" & "011000100000000000000100101100001000000000" & "011000011000000000000100101001000100100000" & "011000010000000000000100100110000010000000" & "011000001000000000000100100011000000100000" & "011000000000000000000100100000000000000000" & "010111111000000000000100011101000000100000" & "010111110000000000000100011010000010000000" & "010111101000000000000100010111000100100000" & "010111100000000000000100010100001000000000" & "010111011000000000000100010001001100100000" & "010111010000000000000100001110010010000000" & "010111001000000000000100001011011000100000" & "010111000000000000000100001000100000000000" & "010110111000000000000100000101101000100000" & "010110110000000000000100000010110010000000" & "010110101000000000000011111111111100100000" & "010110100000000000000011111101001000000000" & "010110011000000000000011111010010100100000" & "010110010000000000000011110111100010000000" & "010110001000000000000011110100110000100000" & "010110000000000000000011110010000000000000" & "010101111000000000000011101111010000100000" & "010101110000000000000011101100100010000000" & "010101101000000000000011101001110100100000" & "010101100000000000000011100111001000000000" & "010101011000000000000011100100011100100000" & "010101010000000000000011100001110010000000" & "010101001000000000000011011111001000100000" & "010101000000000000000011011100100000000000" & "010100111000000000000011011001111000100000" & "010100110000000000000011010111010010000000" & "010100101000000000000011010100101100100000" & "010100100000000000000011010010001000000000" & "010100011000000000000011001111100100100000" & "010100010000000000000011001101000010000000" & "010100001000000000000011001010100000100000" & "010100000000000000000011001000000000000000"
 & "010011111000000000000011000101100000100000" & "010011110000000000000011000011000010000000" & "010011101000000000000011000000100100100000" & "010011100000000000000010111110001000000000" & "010011011000000000000010111011101100100000" & "010011010000000000000010111001010010000000" & "010011001000000000000010110110111000100000" & "010011000000000000000010110100100000000000" & "010010111000000000000010110010001000100000" & "010010110000000000000010101111110010000000" & "010010101000000000000010101101011100100000" & "010010100000000000000010101011001000000000" & "010010011000000000000010101000110100100000" & "010010010000000000000010100110100010000000" & "010010001000000000000010100100010000100000" & "010010000000000000000010100010000000000000" & "010001111000000000000010011111110000100000" & "010001110000000000000010011101100010000000" & "010001101000000000000010011011010100100000" & "010001100000000000000010011001001000000000" & "010001011000000000000010010110111100100000" & "010001010000000000000010010100110010000000" & "010001001000000000000010010010101000100000" & "010001000000000000000010010000100000000000" & "010000111000000000000010001110011000100000" & "010000110000000000000010001100010010000000" & "010000101000000000000010001010001100100000" & "010000100000000000000010001000001000000000" & "010000011000000000000010000110000100100000" & "010000010000000000000010000100000010000000" & "010000001000000000000010000010000000100000" & "010000000000000000000010000000000000000000" & "001111111000000000000001111110000000100000" & "001111110000000000000001111100000010000000" & "001111101000000000000001111010000100100000" & "001111100000000000000001111000001000000000" & "001111011000000000000001110110001100100000" & "001111010000000000000001110100010010000000" & "001111001000000000000001110010011000100000" & "001111000000000000000001110000100000000000" & "001110111000000000000001101110101000100000" & "001110110000000000000001101100110010000000" & "001110101000000000000001101010111100100000" & "001110100000000000000001101001001000000000"
 & "001110011000000000000001100111010100100000" & "001110010000000000000001100101100010000000" & "001110001000000000000001100011110000100000" & "001110000000000000000001100010000000000000" & "001101111000000000000001100000010000100000" & "001101110000000000000001011110100010000000" & "001101101000000000000001011100110100100000" & "001101100000000000000001011011001000000000" & "001101011000000000000001011001011100100000" & "001101010000000000000001010111110010000000" & "001101001000000000000001010110001000100000" & "001101000000000000000001010100100000000000" & "001100111000000000000001010010111000100000" & "001100110000000000000001010001010010000000" & "001100101000000000000001001111101100100000" & "001100100000000000000001001110001000000000" & "001100011000000000000001001100100100100000" & "001100010000000000000001001011000010000000" & "001100001000000000000001001001100000100000" & "001100000000000000000001001000000000000000" & "001011111000000000000001000110100000100000" & "001011110000000000000001000101000010000000" & "001011101000000000000001000011100100100000" & "001011100000000000000001000010001000000000" & "001011011000000000000001000000101100100000" & "001011010000000000000000111111010010000000" & "001011001000000000000000111101111000100000" & "001011000000000000000000111100100000000000" & "001010111000000000000000111011001000100000" & "001010110000000000000000111001110010000000" & "001010101000000000000000111000011100100000" & "001010100000000000000000110111001000000000" & "001010011000000000000000110101110100100000" & "001010010000000000000000110100100010000000" & "001010001000000000000000110011010000100000" & "001010000000000000000000110010000000000000" & "001001111000000000000000110000110000100000" & "001001110000000000000000101111100010000000" & "001001101000000000000000101110010100100000" & "001001100000000000000000101101001000000000" & "001001011000000000000000101011111100100000" & "001001010000000000000000101010110010000000" & "001001001000000000000000101001101000100000" & "001001000000000000000000101000100000000000"
 & "001000111000000000000000100111011000100000" & "001000110000000000000000100110010010000000" & "001000101000000000000000100101001100100000" & "001000100000000000000000100100001000000000" & "001000011000000000000000100011000100100000" & "001000010000000000000000100010000010000000" & "001000001000000000000000100001000000100000" & "001000000000000000000000100000000000000000" & "000111111000000000000000011111000000100000" & "000111110000000000000000011110000010000000" & "000111101000000000000000011101000100100000" & "000111100000000000000000011100001000000000" & "000111011000000000000000011011001100100000" & "000111010000000000000000011010010010000000" & "000111001000000000000000011001011000100000" & "000111000000000000000000011000100000000000" & "000110111000000000000000010111101000100000" & "000110110000000000000000010110110010000000" & "000110101000000000000000010101111100100000" & "000110100000000000000000010101001000000000" & "000110011000000000000000010100010100100000" & "000110010000000000000000010011100010000000" & "000110001000000000000000010010110000100000" & "000110000000000000000000010010000000000000" & "000101111000000000000000010001010000100000" & "000101110000000000000000010000100010000000" & "000101101000000000000000001111110100100000" & "000101100000000000000000001111001000000000" & "000101011000000000000000001110011100100000" & "000101010000000000000000001101110010000000" & "000101001000000000000000001101001000100000" & "000101000000000000000000001100100000000000" & "000100111000000000000000001011111000100000" & "000100110000000000000000001011010010000000" & "000100101000000000000000001010101100100000" & "000100100000000000000000001010001000000000" & "000100011000000000000000001001100100100000" & "000100010000000000000000001001000010000000" & "000100001000000000000000001000100000100000" & "000100000000000000000000001000000000000000" & "000011111000000000000000000111100000100000" & "000011110000000000000000000111000010000000" & "000011101000000000000000000110100100100000" & "000011100000000000000000000110001000000000"
 & "000011011000000000000000000101101100100000" & "000011010000000000000000000101010010000000" & "000011001000000000000000000100111000100000" & "000011000000000000000000000100100000000000" & "000010111000000000000000000100001000100000" & "000010110000000000000000000011110010000000" & "000010101000000000000000000011011100100000" & "000010100000000000000000000011001000000000" & "000010011000000000000000000010110100100000" & "000010010000000000000000000010100010000000" & "000010001000000000000000000010010000100000" & "000010000000000000000000000010000000000000" & "000001111000000000000000000001110000100000" & "000001110000000000000000000001100010000000" & "000001101000000000000000000001010100100000" & "000001100000000000000000000001001000000000" & "000001011000000000000000000000111100100000" & "000001010000000000000000000000110010000000" & "000001001000000000000000000000101000100000" & "000001000000000000000000000000100000000000" & "000000111000000000000000000000011000100000" & "000000110000000000000000000000010010000000" & "000000101000000000000000000000001100100000" & "000000100000000000000000000000001000000000" & "000000011000000000000000000000000100100000" & "000000010000000000000000000000000010000000" & "000000001000000000000000000000000000100000" & "000000000000000000000000000000000000000000");
	table_three_out <= ( "1" & "000000000000000000" & table_three_out_tmp);
	table_three_out_pl <= table_three_dffe12;
	table_three_out_tmp <= wire_table_three_result;
	table_two_data <= ( "111111111011111111001010101011000000010101110111110" & "111111110011111110001010110011000001101011001001011" & "111111101011111101001011000011000100000000001111000" & "111111100011111100001011011011000111010101000000101" & "111111011011111011001011111011001011101001010110001" & "111111010011111010001100100011010000111101000111101" & "111111001011111001001101010011010111010000001100111" & "111111000011111000001110001011011110100010011110001" & "111110111011110111001111001011100110110011110011010" & "111110110011110110010000010011110000000100000100010" & "111110101011110101010001100011111010010011001001001" & "111110100011110100010010111100000101100000111001110" & "111110011011110011010100011100010001101101001110010" & "111110010011110010010110000100011110110111111110101" & "111110001011110001010111110100101101000001000010101" & "111110000011110000011001101100111100001000010010100" & "111101111011101111011011101101001100001101100110001" & "111101110011101110011101110101011101010000110101011" & "111101101011101101100000000101101111010001111000100" & "111101100011101100100010011110000010010000100111010" & "111101011011101011100100111110010110001100111001110" & "111101010011101010100111100110101011000110100111111" & "111101001011101001101010010111000000111101101001110" & "111101000011101000101101001111010111110001110111010" & "111100111011100111110000001111101111100011001000011" & "111100110011100110110011011000001000010001010101000" & "111100101011100101110110101000100001111100010101011" & "111100100011100100111010000000111100100100000001011" & "111100011011100011111101100001011000001000010000111" & "111100010011100011000001001001110100101000111011111" & "111100001011100010000100111010010010000101111010100" & "111100000011100001001000110010110000011111000100101" & "111011111011100000001100110011001111110100010010011" & "111011110011011111010000111011110000000101011011100" & "111011101011011110010101001100010001010010011000001" & "111011100011011101011001100100110011011011000000010" & "111011011011011100011110000101010110011111001011111"
 & "111011010011011011100010101101111010011110110010111" & "111011001011011010100111011110011111011001101101011" & "111011000011011001101100010111000101001111110011010" & "111010111011011000110001010111101100000000111100100" & "111010110011010111110110100000010011101101000001010" & "111010101011010110111011110000111100010011111001010" & "111010100011010110000001001001100101110101011100101" & "111010011011010101000110101010010000010001100011011" & "111010010011010100001100010010111011101000000101100" & "111010001011010011010010000011100111111000111010111" & "111010000011010010010111111100010101000011111011100" & "111001111011010001011101111101000011001000111111100" & "111001110011010000100100000101110010000111111110110" & "111001101011001111101010010110100010000000110001010" & "111001100011001110110000101111010010110011001111000" & "111001011011001101110111010000000100011111010000000" & "111001010011001100111101111000110111000100101100010" & "111001001011001100000100101001101010100011011011101" & "111001000011001011001011100010011110111011010110010" & "111000111011001010010010100011010100001100010100000" & "111000110011001001011001101100001010010110001101000" & "111000101011001000100000111101000001011000111001000" & "111000100011000111101000010101111001010100010000010" & "111000011011000110101111110110110010001000001010100" & "111000010011000101110111011111101011110100100000000" & "111000001011000100111111010000100110011001001000100" & "111000000011000100000111001001100001110101111100001" & "110111111011000011001111001010011110001010110010110" & "110111110011000010010111010011011011010111100100100" & "110111101011000001011111100100011001011100001001010" & "110111100011000000100111111101011000011000011001000" & "110111011010111111110000011110011000001100001011111" & "110111010010111110111001000111011000110111011001101" & "110111001010111110000001111000011010011001111010011" & "110111000010111101001010110001011100110011100110001" & "110110111010111100010011110010100000000100010100110" & "110110110010111011011100111011100100001011111110100"
 & "110110101010111010100110001100101001001010011011000" & "110110100010111001101111100101101110111111100010100" & "110110011010111000111001000110110101101011001100111" & "110110010010111000000010101111111101001101010010001" & "110110001010110111001100100001000101100101101010010" & "110110000010110110010110011010001110110100001101010" & "110101111010110101100000011011011000111000110011001" & "110101110010110100101010100100100011110011010011111" & "110101101010110011110100110101101111100011100111011" & "110101100010110010111111001110111100001001100101101" & "110101011010110010001001110000001001100101000110110" & "110101010010110001010100011001010111110110000010110" & "110101001010110000011111001010100110111100010001011" & "110101000010101111101010000011110110110111101010111" & "110100111010101110110101000101000111101000000111000" & "110100110010101110000000001110011001001101011101111" & "110100101010101101001011011111101011100111100111100" & "110100100010101100010110111000111110110110011011111" & "110100011010101011100010011010010010111001110010111" & "110100010010101010101110000011100111110001100100101" & "110100001010101001111001110100111101011101101001000" & "110100000010101001000101101110010011111101111000000" & "110011111010101000010001101111101011010010001001110" & "110011110010100111011101111001000011011010010110000" & "110011101010100110101010001010011100010110010100111" & "110011100010100101110110100011110110000101111110100" & "110011011010100101000011000101010000101001001010100" & "110011010010100100001111101110101011111111110001010" & "110011001010100011011100100000001000001001101010100" & "110011000010100010101001011001100101000110101110011" & "110010111010100001110110011011000010110110110100101" & "110010110010100001000011100100100001011001110101101" & "110010101010100000010000110110000000101111101001000" & "110010100010011111011110001111100000111000000110111" & "110010011010011110101011110001000001110011000111010" & "110010010010011101111001011010100011100000100010001" & "110010001010011101000111001100000110000000001111100"
 & "110010000010011100010101000101101001010010000111010" & "110001111010011011100011000111001101010110000001100" & "110001110010011010110001010000110010001011110110010" & "110001101010011001111111100010010111110011011101010" & "110001100010011001001101111011111110001100101110110" & "110001011010011000011100011101100101010111100010101" & "110001010010010111101011000111001101010011110001000" & "110001001010010110111001111000110110000001010001101" & "110001000010010110001000110010011111011111111100101" & "110000111010010101010111110100001001101111101001111" & "110000110010010100100110111101110100110000010001101" & "110000101010010011110110001111100000100001101011101" & "110000100010010011000101101001001101000011101111111" & "110000011010010010010101001010111010010110010110100" & "110000010010010001100100110100101000011001010111011" & "110000001010010000110100100110010111001100101010101" & "110000000010010000000100100000000110110000001000000" & "101111111010001111010100100001110111000011100111110" & "101111110010001110100100101011101000000111000001101" & "101111101010001101110100111101011001111010001101110" & "101111100010001101000101010111001100011101000100001" & "101111011010001100010101111000111111101111011100110" & "101111010010001011100110100010110011110001001111100" & "101111001010001010110111010100101000100010010100100" & "101111000010001010001000001110011110000010100011101" & "101110111010001001011001010000010100010001110100111" & "101110110010001000101010011010001011010000000000010" & "101110101010000111111011101100000010111100111101111" & "101110100010000111001101000101111011011000100101100" & "101110011010000110011110100111110100100010101111010" & "101110010010000101110000010001101110011011010011010" & "101110001010000101000010000011101001000010001001001" & "101110000010000100010011111101100100010111001001010" & "101101111010000011100101111111100000011010001011011" & "101101110010000010111000001001011101001011000111100" & "101101101010000010001010011011011010101001110101110" & "101101100010000001011100110101011000110110001110000"
 & "101101011010000000101111010111010111110000001000011" & "101101010010000000000010000001010111010111011100101" & "101101001001111111010100110011010111101100000010111" & "101101000001111110100111101101011000101101110011010" & "101100111001111101111010101111011010011100100101100" & "101100110001111101001101111001011100111000010001110" & "101100101001111100100001001011100000000000101111111" & "101100100001111011110100100101100011110101111000000" & "101100011001111011001000000111101000010111100010001" & "101100010001111010011011110001101101100101100110001" & "101100001001111001101111100011110011011111111100000" & "101100000001111001000011011101111010000110011011111" & "101011111001111000010111100000000001011000111101100" & "101011110001110111101011101010001001010111011001001" & "101011101001110110111111111100010010000001100110101" & "101011100001110110010100010110011011010111011101111" & "101011011001110101101000111000100101011000110111000" & "101011010001110100111101100010110000000101101010000" & "101011001001110100010010010100111011011101101110111" & "101011000001110011100111001111000111100000111101100" & "101010111001110010111100010001010100001111001110000" & "101010110001110010010001011011100001101000011000010" & "101010101001110001100110101101101111101100010100010" & "101010100001110000111100000111111110011010111010001" & "101010011001110000010001101010001101110100000001101" & "101010010001101111100111010100011101110111100011000" & "101010001001101110111101000110101110100101010110000" & "101010000001101110010011000000111111111101010010111" & "101001111001101101101001000011010001111111010001011" & "101001110001101100111111001101100100101011001001101" & "101001101001101100010101011111111000000000110011100" & "101001100001101011101011111010001100000000000111010" & "101001011001101011000010011100100000101000111100100" & "101001010001101010011001000110110101111011001011100" & "101001001001101001101111111001001011110110101100001" & "101001000001101001000110110011100010011011010110100" & "101000111001101000011101110101111001101001000010011"
 & "101000110001100111110101000000010001011111101000000" & "101000101001100111001100010010101001111110111111010" & "101000100001100110100011101101000011000111000000000" & "101000011001100101111011001111011100110111100010011" & "101000010001100101010010111001110111010000011110011" & "101000001001100100101010101100010010010001101100000" & "101000000001100100000010100110101101111011000011010" & "100111111001100011011010101001001010001100011011111" & "100111110001100010110010110011100111000101101110010" & "100111101001100010001011000110000100100110110010000" & "100111100001100001100011100000100010101111011111011" & "100111011001100000111100000011000001011111101110010" & "100111010001100000010100101101100000110111010110101" & "100111001001011111101101100000000000110110010000101" & "100111000001011111000110011010100001011100010100000" & "100110111001011110011111011101000010101001011000111" & "100110110001011101111000100111100100011101010111010" & "100110101001011101010001111010000110111000000111000" & "100110100001011100101011010100101001111001100000011" & "100110011001011100000100110111001101100001011011001" & "100110010001011011011110100001110001101111101111010" & "100110001001011010111000010100010110100100010100111" & "100110000001011010010010001110111011111111000011111" & "100101111001011001101100010001100001111111110100010" & "100101110001011001000110011100001000100110011110001" & "100101101001011000100000101110101111110010111001011" & "100101100001010111111011001001010111100100111110000" & "100101011001010111010101101011111111111100100100000" & "100101010001010110110000010110101000111001100011010" & "100101001001010110001011001001010010011011110100000" & "100101000001010101100110000011111100100011001110001" & "100100111001010101000001000110100111001111101001100" & "100100110001010100011100010001010010100000111110001" & "100100101001010011110111100011111110010111000100010" & "100100100001010011010010111110101010110001110011100" & "100100011001010010101110100001010111110001000100010" & "100100010001010010001010001100000101010100101110001"
 & "100100001001010001100101111110110011011100101001011" & "100100000001010001000001111001100010001000101101111" & "100011111001010000011101111100010001011000110011101" & "100011110001001111111010000111000001001100110010101" & "100011101001001111010110011001110001100100100010111" & "100011100001001110110010110100100010011111111100011" & "100011011001001110001111010111010011111110110111001" & "100011010001001101101100000010000110000001001011001" & "100011001001001101001000110100111000100110110000010" & "100011000001001100100101101111101011101111011110110" & "100010111001001100000010110010011111011011001110010" & "100010110001001011011111111101010011101001110111000" & "100010101001001010111101010000001000011011010001000" & "100010100001001010011010101010111101101111010100001" & "100010011001001001111000001101110011100101111000011" & "100010010001001001010101111000101001111110110101111" & "100010001001001000110011101011100000111010000100011" & "100010000001001000010001100110011000010111011100001" & "100001111001000111101111101001010000010110110101000" & "100001110001000111001101110100001000111000000111000" & "100001101001000110101100000111000001111011001010000" & "100001100001000110001010100001111011011111110110010" & "100001011001000101101001000100110101100110000011100" & "100001010001000101000111101111110000001101101001111" & "100001001001000100100110100010101011010110100001011" & "100001000001000100000101011101100111000000100001111" & "100000111001000011100100100000100011001011100011100" & "100000110001000011000011101011011111110111011110001" & "100000101001000010100010111110011101000100001001110" & "100000100001000010000010011001011010110001011110100" & "100000011001000001100001111100011000111111010100010" & "100000010001000001000001100111010111101101100011000" & "100000001001000000100001011010010110111100000010111" & "100000000001000000000001010101010110101010101011101" & "011111111000111111100001011000010110111001010101100" & "011111110000111111000001100011010111100111111000010" & "011111101000111110100001110110011000110110001100001"
 & "011111100000111110000010010001011010100100001000111" & "011111011000111101100010110100011100110001100110101" & "011111010000111101000011011111011111011110011101010" & "011111001000111100100100010010100010101010100100111" & "011111000000111100000101001101100110010101110101100" & "011110111000111011100110010000101010100000000111000" & "011110110000111011000111011011101111001001010001100" & "011110101000111010101000101110110100010001001100111" & "011110100000111010001010001001111001110111110001010" & "011110011000111001101011101100111111111100110110011" & "011110010000111001001101011000000110100000010100100" & "011110001000111000101111001011001101100010000011100" & "011110000000111000010001000110010101000001111011100" & "011101111000110111110011001001011100111111110100010" & "011101110000110111010101010100100101011011100101111" & "011101101000110110110111100111101110010101001000011" & "011101100000110110011010000010110111101100010011110" & "011101011000110101111100100110000001100001000000000" & "011101010000110101011111010001001011110011000101000" & "011101001000110101000010000100010110100010011011000" & "011101000000110100100100111111100001101110111001101" & "011100111000110100001000000010101101011000011001010" & "011100110000110011101011001101111001011110110001101" & "011100101000110011001110100001000110000001111010110" & "011100100000110010110001111100010011000001101100110" & "011100011000110010010101011111100000011101111111100" & "011100010000110001111001001010101110010110101011000" & "011100001000110001011100111101111100101011100111011" & "011100000000110001000000111001001011011100101100100" & "011011111000110000100100111100011010101001110010011" & "011011110000110000001001000111101010010010110001000" & "011011101000101111101101011010111010010111100000011" & "011011100000101111010001110110001010110111111000100" & "011011011000101110110110011001011011110011110001011" & "011011010000101110011011000100101101001011000011000" & "011011001000101101111111110111111110111101100101010" & "011011000000101101100100110011010001001011010000011"
 & "011010111000101101001001110110100011110011111100001" & "011010110000101100101111000001110110110111100000100" & "011010101000101100010100010101001010010101110101101" & "011010100000101011111001110000011110001110110011100" & "011010011000101011011111010011110010100010010010001" & "011010010000101011000100111111000111010000001001010" & "011010001000101010101010110010011100011000010001001" & "011010000000101010010000101101110001111010100001110" & "011001111000101001110110110001000111110110110011000" & "011001110000101001011100111100011110001100111100111" & "011001101000101001000011001111110100111100110111011" & "011001100000101000101001101011001100000110011010100" & "011001011000101000010000001110100011101001011110010" & "011001010000100111110110111001111011100101111010110" & "011001001000100111011101101101010011111011100111110" & "011001000000100111000100101000101100101010011101011" & "011000111000100110101011101100000101110010010011110" & "011000110000100110010010110111011111010011000010101" & "011000101000100101111010001010111001001100100010000" & "011000100000100101100001100110010011011110101010001" & "011000011000100101001001001001101110001001010010110" & "011000010000100100110000110101001001001100010100000" & "011000001000100100011000101000100100100111100101111" & "011000000000100100000000100100000000011011000000010" & "010111111000100011101000100111011100100110011011001" & "010111110000100011010000110010111001001001101110101" & "010111101000100010111001000110010110000100110010101" & "010111100000100010100001100001110011010111011111010" & "010111011000100010001010000101010001000001101100011" & "010111010000100001110010110000101111000011010010001" & "010111001000100001011011100100001101011100001000010" & "010111000000100001000100011111101100001100000111000" & "010110111000100000101101100011001011010011000110010" & "010110110000100000010110101110101010110000111110000" & "010110101000100000000000000010001010100101100110010" & "010110100000011111101001011101101010110000110111000" & "010110011000011111010011000001001011010010101000010"
 & "010110010000011110111100101100101100001010110010000" & "010110001000011110100110100000001101011001001100001" & "010110000000011110010000011011101110111101101110111" & "010101111000011101111010011111010000111000010010000" & "010101110000011101100100101010110011001000101101101" & "010101101000011101001110111110010101101110111001110" & "010101100000011100111001011001111000101010101110010" & "010101011000011100100011111101011011111100000011011" & "010101010000011100001110101000111111100010110000110" & "010101001000011011111001011100100011011110101110101" & "010101000000011011100100011000000111101111110101000" & "010100111000011011001111011011101100010101111011110" & "010100110000011010111010100111010001010000111010111" & "010100101000011010100101111010110110100000101010100" & "010100100000011010010001010110011100000101000010101" & "010100011000011001111100111010000001111101111011000" & "010100010000011001101000100101101000001011001011111" & "010100001000011001010100011001001110101100101101001" & "010100000000011001000000010100110101100010010110110" & "010011111000011000101100011000011100101100000000110" & "010011110000011000011000100100000100001001100011001" & "010011101000011000000100110111101011111010110101111" & "010011100000010111110001010011010011111111110001001" & "010011011000010111011101110110111100011000001100101" & "010011010000010111001010100010100101000100000000100" & "010011001000010110110111010110001110000011000100111" & "010011000000010110100100010001110111010101010001100" & "010010111000010110010001010101100000111010011110011" & "010010110000010101111110100001001010110010100011110" & "010010101000010101101011110100110100111101011001011" & "010010100000010101011001010000011111011010110111011" & "010010011000010101000110110100001010001010110101110" & "010010010000010100110100011111110101001101001100011" & "010010001000010100100010010011100000100001110011011" & "010010000000010100010000001111001100001000100010110" & "010001111000010011111110010010111000000001010010011" & "010001110000010011101100011110100100001011111010011"
 & "010001101000010011011010110010010000101000010010101" & "010001100000010011001001001101111101010110010011001" & "010001011000010010110111110001101010010101110100000" & "010001010000010010100110011101010111100110101101001" & "010001001000010010010101010001000101001000110110101" & "010001000000010010000100001100110010111100001000011" & "010000111000010001110011010000100001000000011010011" & "010000110000010001100010011100001111010101100100101" & "010000101000010001010001101111111101111011011111001" & "010000100000010001000001001011101100110010000010000" & "010000011000010000110000101111011011111001000101001" & "010000010000010000100000011011001011010000100000100" & "010000001000010000010000001110111010111000001100001" & "010000000000010000000000001010101010110000000000000" & "001111111000001111110000001110011010110111110100001" & "001111110000001111100000011010001011001111100000100" & "001111101000001111010000101101111011110110111101001" & "001111100000001111000001001001101100101110000001111" & "001111011000001110110001101101011101110100100111000" & "001111010000001110100010011001001111001010100100011" & "001111001000001110010011001101000000101111110001111" & "001111000000001110000100001000110010100100000111101" & "001110111000001101110101001100100100100111011101101" & "001110110000001101100110011000010110111001101011111" & "001110101000001101010111101100001001011010101010010" & "001110100000001101001001000111111100001010010000111" & "001110011000001100111010101011101111001000010111110" & "001110010000001100101100010111100010010100110110110" & "001110001000001100011110001011010101101111100110000" & "001110000000001100010000000111001001011000011101011" & "001101111000001100000010001010111101001111010101000" & "001101110000001011110100010110110001010100000100110" & "001101101000001011100110101010100101100110100100110" & "001101100000001011011001000110011010000110101101000" & "001101011000001011001011101010001110110100010101010" & "001101010000001010111110010110000011101111010101111" & "001101001000001010110001001001111000110111100110100"
 & "001101000000001010100100000101101110001100111111011" & "001100111000001010010111001001100011101111011000011" & "001100110000001010001010010101011001011110101001101" & "001100101000001001111101101001001111011010101010111" & "001100100000001001110001000101000101100011010100011" & "001100011000001001100100101000111011111000011110001" & "001100010000001001011000010100110010011001111111111" & "001100001000001001001100001000101001000111110001111" & "001100000000001001000000000100100000000001101100000" & "001011111000001000110100001000010111000111100110001" & "001011110000001000101000010100001110011001011000100" & "001011101000001000011100101000000101110110111011001" & "001011100000001000010001000011111101100000000101110" & "001011011000001000000101100111110101010100110000100" & "001011010000000111111010010011101101010100110011011" & "001011001000000111101111000111100101100000000110011" & "001011000000000111100100000011011101110110100001100" & "001010111000000111011001000111010110010111111100110" & "001010110000000111001110010011001111000100010000001" & "001010101000000111000011100111000111111011010011101" & "001010100000000110111001000011000000111100111111010" & "001010011000000110101110100110111010001001001011000" & "001010010000000110100100010010110011011111101110110" & "001010001000000110011010000110101101000000100010101" & "001010000000000110010000000010100110101011011110110" & "001001111000000110000110000110100000100000011010110" & "001001110000000101111100010010011010011111001111000" & "001001101000000101110010100110010100100111110011010" & "001001100000000101101001000010001110111001111111110" & "001001011000000101011111100110001001010101101100001" & "001001010000000101010110010010000011111010110000110" & "001001001000000101001101000101111110101001000101011" & "001001000000000101000100000001111001100000100010001" & "001000111000000100111011000101110100100000111110111" & "001000110000000100110010010001101111101010010011110" & "001000101000000100101001100101101010111100011000110" & "001000100000000100100001000001100110010111000101110"
 & "001000011000000100011000100101100001111010010010111" & "001000010000000100010000010001011101100101111000001" & "001000001000000100001000000101011001011001101101010" & "001000000000000100000000000001010101010101101010101" & "000111111000000011111000000101010001011001101000000" & "000111110000000011110000010001001101100101011101011" & "000111101000000011101000100101001001111001000010111" & "000111100000000011100001000001000110010100010000011" & "000111011000000011011001100101000010110110111110000" & "000111010000000011010010010000111111100001000011101" & "000111001000000011001011000100111100010010011001011" & "000111000000000011000100000000111001001010110111001" & "000110111000000010111101000100110110001010010100111" & "000110110000000010110110010000110011010000101010110" & "000110101000000010101111100100110000011101110000101" & "000110100000000010101001000000101101110001011110101" & "000110011000000010100010100100101011001011101100100" & "000110010000000010011100010000101000101100010010100" & "000110001000000010010110000100100110010011001000101" & "000110000000000010010000000000100100000000000110101" & "000101111000000010001010000100100001110011000100110" & "000101110000000010000100010000011111101011111011000" & "000101101000000001111110100100011101101010100001001" & "000101100000000001111001000000011011101110101111011" & "000101011000000001110011100100011001111000011101101" & "000101010000000001101110010000011000000111100011111" & "000101001000000001101001000100010110011011111010010" & "000101000000000001100100000000010100110101011000100" & "000100111000000001011111000100010011010011110110111" & "000100110000000001011010010000010001110111001101010" & "000100101000000001010101100100010000011111010011101" & "000100100000000001010001000000001111001100000010001" & "000100011000000001001100100100001101111101010000100" & "000100010000000001001000010000001100110010110111000" & "000100001000000001000100000100001011101100101101100" & "000100000000000001000000000000001010101010101011111" & "000011111000000000111100000100001001101100101010100"
 & "000011110000000000111000010000001000110010100001000" & "000011101000000000110100100100000111111100000111100" & "000011100000000000110001000000000111001001010110000" & "000011011000000000101101100100000110011010000100101" & "000011010000000000101010010000000101101110001011001" & "000011001000000000100111000100000101000101100001110" & "000011000000000000100100000000000100100000000000011" & "000010111000000000100001000100000011111101011111000" & "000010110000000000011110010000000011011101110101101" & "000010101000000000011011100100000011000000111100001" & "000010100000000000011001000000000010100110101010110" & "000010011000000000010110100100000010001110111001011" & "000010010000000000010100010000000001111001100000001" & "000010001000000000010010000100000001100110010110110" & "000010000000000000010000000000000001010101010101011" & "000001111000000000001110000100000001000110010100000" & "000001110000000000001100010000000000111001001010101" & "000001101000000000001010100100000000101101110001010" & "000001100000000000001001000000000000100100000000000" & "000001011000000000000111100100000000011011101110101" & "000001010000000000000110010000000000010100110101010" & "000001001000000000000101000100000000001111001100000" & "000001000000000000000100000000000000001010101010101" & "000000111000000000000011000100000000000111001001010" & "000000110000000000000010010000000000000100100000000" & "000000101000000000000001100100000000000010100110101" & "000000100000000000000001000000000000000001010101010" & "000000011000000000000000100100000000000000100011111" & "000000010000000000000000010000000000000000001010101" & "000000001000000000000000000100000000000000000001010" & "000000000000000000000000000000000000000000000000000");
	table_two_out <= ( "1" & "000000000" & table_two_out_tmp);
	table_two_out_pl <= table_two_dffe12;
	table_two_out_tmp <= wire_table_two_result;
	tbl1_compare_wi <= wire_tbl1_compare_ageb;
	tbl1_compare_wo <= tbl1_compare_dffe11_10_pipes9;
	tbl1_tbl2_prod_wi <= wire_tbl1_tbl2_prod_result(121 DOWNTO 62);
	tbl1_tbl2_prod_wo <= tbl1_tbl2_prod_wi;
	tbl3_taylor_prod_wi <= wire_tbl3_taylor_prod_result(119 DOWNTO 60);
	tbl3_taylor_prod_wo <= tbl3_taylor_prod_wi;
	underflow_compare_val_w <= "00000111010";
	underflow_w <= (((((result_underflow_w OR barrel_shifter_underflow) OR wire_sign_dffe_w_lg_q3430w(0)) AND wire_w_lg_input_is_zero_wo3426w(0)) AND wire_w_lg_input_is_infinity_wo3425w(0)) AND wire_w_lg_input_is_nan_wo3424w(0));
	x_fixed <= wire_rbarrel_shift_result;
	xf <= wire_xf_muxa_dataout;
	xf_pl <= xf_pl_dffe12;
	xf_pre <= wire_x_fixed_minus_xiln2_result;
	xf_pre_2_wi <= xf_pre_wo;
	xf_pre_2_wo <= xf_pre_2_dffe10;
	xf_pre_wi <= xf_pre;
	xf_pre_wo <= xf_pre_dffe9;
	xi_exp_value <= xi_prod_wo(24 DOWNTO 14);
	xi_exp_value_wi <= xi_exp_value;
	xi_exp_value_wo <= xi_exp_value_dffe4;
	xi_ln2_prod_wi <= wire_xi_ln2_prod_result;
	xi_ln2_prod_wo <= xi_ln2_prod_dffe7;
	xi_prod_wi <= wire_xi_prod_result;
	xi_prod_wo <= xi_prod_dffe3;
	wire_w_data_range93w(0) <= data(10);
	wire_w_data_range96w(0) <= data(11);
	wire_w_data_range99w(0) <= data(12);
	wire_w_data_range102w(0) <= data(13);
	wire_w_data_range105w(0) <= data(14);
	wire_w_data_range108w(0) <= data(15);
	wire_w_data_range111w(0) <= data(16);
	wire_w_data_range114w(0) <= data(17);
	wire_w_data_range117w(0) <= data(18);
	wire_w_data_range120w(0) <= data(19);
	wire_w_data_range66w(0) <= data(1);
	wire_w_data_range123w(0) <= data(20);
	wire_w_data_range126w(0) <= data(21);
	wire_w_data_range129w(0) <= data(22);
	wire_w_data_range132w(0) <= data(23);
	wire_w_data_range135w(0) <= data(24);
	wire_w_data_range138w(0) <= data(25);
	wire_w_data_range141w(0) <= data(26);
	wire_w_data_range144w(0) <= data(27);
	wire_w_data_range147w(0) <= data(28);
	wire_w_data_range150w(0) <= data(29);
	wire_w_data_range69w(0) <= data(2);
	wire_w_data_range153w(0) <= data(30);
	wire_w_data_range156w(0) <= data(31);
	wire_w_data_range159w(0) <= data(32);
	wire_w_data_range162w(0) <= data(33);
	wire_w_data_range165w(0) <= data(34);
	wire_w_data_range168w(0) <= data(35);
	wire_w_data_range171w(0) <= data(36);
	wire_w_data_range174w(0) <= data(37);
	wire_w_data_range177w(0) <= data(38);
	wire_w_data_range180w(0) <= data(39);
	wire_w_data_range72w(0) <= data(3);
	wire_w_data_range183w(0) <= data(40);
	wire_w_data_range186w(0) <= data(41);
	wire_w_data_range189w(0) <= data(42);
	wire_w_data_range192w(0) <= data(43);
	wire_w_data_range195w(0) <= data(44);
	wire_w_data_range198w(0) <= data(45);
	wire_w_data_range201w(0) <= data(46);
	wire_w_data_range204w(0) <= data(47);
	wire_w_data_range207w(0) <= data(48);
	wire_w_data_range210w(0) <= data(49);
	wire_w_data_range75w(0) <= data(4);
	wire_w_data_range213w(0) <= data(50);
	wire_w_data_range216w(0) <= data(51);
	wire_w_data_range10w(0) <= data(53);
	wire_w_data_range13w(0) <= data(54);
	wire_w_data_range16w(0) <= data(55);
	wire_w_data_range19w(0) <= data(56);
	wire_w_data_range22w(0) <= data(57);
	wire_w_data_range25w(0) <= data(58);
	wire_w_data_range28w(0) <= data(59);
	wire_w_data_range78w(0) <= data(5);
	wire_w_data_range31w(0) <= data(60);
	wire_w_data_range34w(0) <= data(61);
	wire_w_data_range37w(0) <= data(62);
	wire_w_data_range81w(0) <= data(6);
	wire_w_data_range84w(0) <= data(7);
	wire_w_data_range87w(0) <= data(8);
	wire_w_data_range90w(0) <= data(9);
	wire_w_exp_data_all_one_w_range41w(0) <= exp_data_all_one_w(0);
	wire_w_exp_data_all_one_w_range62w(0) <= exp_data_all_one_w(10);
	wire_w_exp_data_all_one_w_range44w(0) <= exp_data_all_one_w(1);
	wire_w_exp_data_all_one_w_range46w(0) <= exp_data_all_one_w(2);
	wire_w_exp_data_all_one_w_range48w(0) <= exp_data_all_one_w(3);
	wire_w_exp_data_all_one_w_range50w(0) <= exp_data_all_one_w(4);
	wire_w_exp_data_all_one_w_range52w(0) <= exp_data_all_one_w(5);
	wire_w_exp_data_all_one_w_range54w(0) <= exp_data_all_one_w(6);
	wire_w_exp_data_all_one_w_range56w(0) <= exp_data_all_one_w(7);
	wire_w_exp_data_all_one_w_range58w(0) <= exp_data_all_one_w(8);
	wire_w_exp_data_all_one_w_range60w(0) <= exp_data_all_one_w(9);
	wire_w_exp_data_not_zero_w_range8w(0) <= exp_data_not_zero_w(0);
	wire_w_exp_data_not_zero_w_range12w(0) <= exp_data_not_zero_w(1);
	wire_w_exp_data_not_zero_w_range15w(0) <= exp_data_not_zero_w(2);
	wire_w_exp_data_not_zero_w_range18w(0) <= exp_data_not_zero_w(3);
	wire_w_exp_data_not_zero_w_range21w(0) <= exp_data_not_zero_w(4);
	wire_w_exp_data_not_zero_w_range24w(0) <= exp_data_not_zero_w(5);
	wire_w_exp_data_not_zero_w_range27w(0) <= exp_data_not_zero_w(6);
	wire_w_exp_data_not_zero_w_range30w(0) <= exp_data_not_zero_w(7);
	wire_w_exp_data_not_zero_w_range33w(0) <= exp_data_not_zero_w(8);
	wire_w_exp_data_not_zero_w_range36w(0) <= exp_data_not_zero_w(9);
	wire_w_exp_out_all_one_w_range3628w(0) <= exp_out_all_one_w(0);
	wire_w_exp_out_all_one_w_range3634w(0) <= exp_out_all_one_w(1);
	wire_w_exp_out_all_one_w_range3639w(0) <= exp_out_all_one_w(2);
	wire_w_exp_out_all_one_w_range3644w(0) <= exp_out_all_one_w(3);
	wire_w_exp_out_all_one_w_range3649w(0) <= exp_out_all_one_w(4);
	wire_w_exp_out_all_one_w_range3654w(0) <= exp_out_all_one_w(5);
	wire_w_exp_out_all_one_w_range3659w(0) <= exp_out_all_one_w(6);
	wire_w_exp_out_all_one_w_range3664w(0) <= exp_out_all_one_w(7);
	wire_w_exp_out_all_one_w_range3669w(0) <= exp_out_all_one_w(8);
	wire_w_exp_out_all_one_w_range3674w(0) <= exp_out_all_one_w(9);
	wire_w_exp_out_not_zero_w_range3630w(0) <= exp_out_not_zero_w(0);
	wire_w_exp_out_not_zero_w_range3636w(0) <= exp_out_not_zero_w(1);
	wire_w_exp_out_not_zero_w_range3641w(0) <= exp_out_not_zero_w(2);
	wire_w_exp_out_not_zero_w_range3646w(0) <= exp_out_not_zero_w(3);
	wire_w_exp_out_not_zero_w_range3651w(0) <= exp_out_not_zero_w(4);
	wire_w_exp_out_not_zero_w_range3656w(0) <= exp_out_not_zero_w(5);
	wire_w_exp_out_not_zero_w_range3661w(0) <= exp_out_not_zero_w(6);
	wire_w_exp_out_not_zero_w_range3666w(0) <= exp_out_not_zero_w(7);
	wire_w_exp_out_not_zero_w_range3671w(0) <= exp_out_not_zero_w(8);
	wire_w_exp_out_not_zero_w_range3676w(0) <= exp_out_not_zero_w(9);
	wire_w_exp_result_w_range3677w(0) <= exp_result_w(10);
	wire_w_exp_result_w_range3632w(0) <= exp_result_w(1);
	wire_w_exp_result_w_range3637w(0) <= exp_result_w(2);
	wire_w_exp_result_w_range3642w(0) <= exp_result_w(3);
	wire_w_exp_result_w_range3647w(0) <= exp_result_w(4);
	wire_w_exp_result_w_range3652w(0) <= exp_result_w(5);
	wire_w_exp_result_w_range3657w(0) <= exp_result_w(6);
	wire_w_exp_result_w_range3662w(0) <= exp_result_w(7);
	wire_w_exp_result_w_range3667w(0) <= exp_result_w(8);
	wire_w_exp_result_w_range3672w(0) <= exp_result_w(9);
	wire_w_exp_value_wo_range234w <= exp_value_wo(10 DOWNTO 0);
	wire_w_exp_value_wo_range233w(0) <= exp_value_wo(11);
	wire_w_exp_value_wo_range231w <= exp_value_wo(6 DOWNTO 0);
	wire_w_man_data_not_zero_w_range64w(0) <= man_data_not_zero_w(0);
	wire_w_man_data_not_zero_w_range95w(0) <= man_data_not_zero_w(10);
	wire_w_man_data_not_zero_w_range98w(0) <= man_data_not_zero_w(11);
	wire_w_man_data_not_zero_w_range101w(0) <= man_data_not_zero_w(12);
	wire_w_man_data_not_zero_w_range104w(0) <= man_data_not_zero_w(13);
	wire_w_man_data_not_zero_w_range107w(0) <= man_data_not_zero_w(14);
	wire_w_man_data_not_zero_w_range110w(0) <= man_data_not_zero_w(15);
	wire_w_man_data_not_zero_w_range113w(0) <= man_data_not_zero_w(16);
	wire_w_man_data_not_zero_w_range116w(0) <= man_data_not_zero_w(17);
	wire_w_man_data_not_zero_w_range119w(0) <= man_data_not_zero_w(18);
	wire_w_man_data_not_zero_w_range122w(0) <= man_data_not_zero_w(19);
	wire_w_man_data_not_zero_w_range68w(0) <= man_data_not_zero_w(1);
	wire_w_man_data_not_zero_w_range125w(0) <= man_data_not_zero_w(20);
	wire_w_man_data_not_zero_w_range128w(0) <= man_data_not_zero_w(21);
	wire_w_man_data_not_zero_w_range131w(0) <= man_data_not_zero_w(22);
	wire_w_man_data_not_zero_w_range134w(0) <= man_data_not_zero_w(23);
	wire_w_man_data_not_zero_w_range137w(0) <= man_data_not_zero_w(24);
	wire_w_man_data_not_zero_w_range140w(0) <= man_data_not_zero_w(25);
	wire_w_man_data_not_zero_w_range143w(0) <= man_data_not_zero_w(26);
	wire_w_man_data_not_zero_w_range146w(0) <= man_data_not_zero_w(27);
	wire_w_man_data_not_zero_w_range149w(0) <= man_data_not_zero_w(28);
	wire_w_man_data_not_zero_w_range152w(0) <= man_data_not_zero_w(29);
	wire_w_man_data_not_zero_w_range71w(0) <= man_data_not_zero_w(2);
	wire_w_man_data_not_zero_w_range155w(0) <= man_data_not_zero_w(30);
	wire_w_man_data_not_zero_w_range158w(0) <= man_data_not_zero_w(31);
	wire_w_man_data_not_zero_w_range161w(0) <= man_data_not_zero_w(32);
	wire_w_man_data_not_zero_w_range164w(0) <= man_data_not_zero_w(33);
	wire_w_man_data_not_zero_w_range167w(0) <= man_data_not_zero_w(34);
	wire_w_man_data_not_zero_w_range170w(0) <= man_data_not_zero_w(35);
	wire_w_man_data_not_zero_w_range173w(0) <= man_data_not_zero_w(36);
	wire_w_man_data_not_zero_w_range176w(0) <= man_data_not_zero_w(37);
	wire_w_man_data_not_zero_w_range179w(0) <= man_data_not_zero_w(38);
	wire_w_man_data_not_zero_w_range182w(0) <= man_data_not_zero_w(39);
	wire_w_man_data_not_zero_w_range74w(0) <= man_data_not_zero_w(3);
	wire_w_man_data_not_zero_w_range185w(0) <= man_data_not_zero_w(40);
	wire_w_man_data_not_zero_w_range188w(0) <= man_data_not_zero_w(41);
	wire_w_man_data_not_zero_w_range191w(0) <= man_data_not_zero_w(42);
	wire_w_man_data_not_zero_w_range194w(0) <= man_data_not_zero_w(43);
	wire_w_man_data_not_zero_w_range197w(0) <= man_data_not_zero_w(44);
	wire_w_man_data_not_zero_w_range200w(0) <= man_data_not_zero_w(45);
	wire_w_man_data_not_zero_w_range203w(0) <= man_data_not_zero_w(46);
	wire_w_man_data_not_zero_w_range206w(0) <= man_data_not_zero_w(47);
	wire_w_man_data_not_zero_w_range209w(0) <= man_data_not_zero_w(48);
	wire_w_man_data_not_zero_w_range212w(0) <= man_data_not_zero_w(49);
	wire_w_man_data_not_zero_w_range77w(0) <= man_data_not_zero_w(4);
	wire_w_man_data_not_zero_w_range215w(0) <= man_data_not_zero_w(50);
	wire_w_man_data_not_zero_w_range218w(0) <= man_data_not_zero_w(51);
	wire_w_man_data_not_zero_w_range80w(0) <= man_data_not_zero_w(5);
	wire_w_man_data_not_zero_w_range83w(0) <= man_data_not_zero_w(6);
	wire_w_man_data_not_zero_w_range86w(0) <= man_data_not_zero_w(7);
	wire_w_man_data_not_zero_w_range89w(0) <= man_data_not_zero_w(8);
	wire_w_man_data_not_zero_w_range92w(0) <= man_data_not_zero_w(9);
	wire_w_man_prod_result_range3406w(0) <= man_prod_result(58);
	wire_w_man_prod_result_range3403w(0) <= man_prod_result(59);
	wire_w_man_prod_result_range3400w(0) <= man_prod_result(60);
	wire_w_man_prod_result_range3397w(0) <= man_prod_result(61);
	wire_w_man_prod_wo_range3384w(0) <= man_prod_wo(117);
	wire_w_man_result_all_ones_range3445w(0) <= man_result_all_ones(0);
	wire_w_man_result_all_ones_range3476w(0) <= man_result_all_ones(10);
	wire_w_man_result_all_ones_range3479w(0) <= man_result_all_ones(11);
	wire_w_man_result_all_ones_range3482w(0) <= man_result_all_ones(12);
	wire_w_man_result_all_ones_range3485w(0) <= man_result_all_ones(13);
	wire_w_man_result_all_ones_range3488w(0) <= man_result_all_ones(14);
	wire_w_man_result_all_ones_range3491w(0) <= man_result_all_ones(15);
	wire_w_man_result_all_ones_range3494w(0) <= man_result_all_ones(16);
	wire_w_man_result_all_ones_range3497w(0) <= man_result_all_ones(17);
	wire_w_man_result_all_ones_range3500w(0) <= man_result_all_ones(18);
	wire_w_man_result_all_ones_range3503w(0) <= man_result_all_ones(19);
	wire_w_man_result_all_ones_range3449w(0) <= man_result_all_ones(1);
	wire_w_man_result_all_ones_range3506w(0) <= man_result_all_ones(20);
	wire_w_man_result_all_ones_range3509w(0) <= man_result_all_ones(21);
	wire_w_man_result_all_ones_range3512w(0) <= man_result_all_ones(22);
	wire_w_man_result_all_ones_range3515w(0) <= man_result_all_ones(23);
	wire_w_man_result_all_ones_range3518w(0) <= man_result_all_ones(24);
	wire_w_man_result_all_ones_range3521w(0) <= man_result_all_ones(25);
	wire_w_man_result_all_ones_range3524w(0) <= man_result_all_ones(26);
	wire_w_man_result_all_ones_range3527w(0) <= man_result_all_ones(27);
	wire_w_man_result_all_ones_range3530w(0) <= man_result_all_ones(28);
	wire_w_man_result_all_ones_range3533w(0) <= man_result_all_ones(29);
	wire_w_man_result_all_ones_range3452w(0) <= man_result_all_ones(2);
	wire_w_man_result_all_ones_range3536w(0) <= man_result_all_ones(30);
	wire_w_man_result_all_ones_range3539w(0) <= man_result_all_ones(31);
	wire_w_man_result_all_ones_range3542w(0) <= man_result_all_ones(32);
	wire_w_man_result_all_ones_range3545w(0) <= man_result_all_ones(33);
	wire_w_man_result_all_ones_range3548w(0) <= man_result_all_ones(34);
	wire_w_man_result_all_ones_range3551w(0) <= man_result_all_ones(35);
	wire_w_man_result_all_ones_range3554w(0) <= man_result_all_ones(36);
	wire_w_man_result_all_ones_range3557w(0) <= man_result_all_ones(37);
	wire_w_man_result_all_ones_range3560w(0) <= man_result_all_ones(38);
	wire_w_man_result_all_ones_range3563w(0) <= man_result_all_ones(39);
	wire_w_man_result_all_ones_range3455w(0) <= man_result_all_ones(3);
	wire_w_man_result_all_ones_range3566w(0) <= man_result_all_ones(40);
	wire_w_man_result_all_ones_range3569w(0) <= man_result_all_ones(41);
	wire_w_man_result_all_ones_range3572w(0) <= man_result_all_ones(42);
	wire_w_man_result_all_ones_range3575w(0) <= man_result_all_ones(43);
	wire_w_man_result_all_ones_range3578w(0) <= man_result_all_ones(44);
	wire_w_man_result_all_ones_range3581w(0) <= man_result_all_ones(45);
	wire_w_man_result_all_ones_range3584w(0) <= man_result_all_ones(46);
	wire_w_man_result_all_ones_range3587w(0) <= man_result_all_ones(47);
	wire_w_man_result_all_ones_range3590w(0) <= man_result_all_ones(48);
	wire_w_man_result_all_ones_range3593w(0) <= man_result_all_ones(49);
	wire_w_man_result_all_ones_range3458w(0) <= man_result_all_ones(4);
	wire_w_man_result_all_ones_range3596w(0) <= man_result_all_ones(50);
	wire_w_man_result_all_ones_range3461w(0) <= man_result_all_ones(5);
	wire_w_man_result_all_ones_range3464w(0) <= man_result_all_ones(6);
	wire_w_man_result_all_ones_range3467w(0) <= man_result_all_ones(7);
	wire_w_man_result_all_ones_range3470w(0) <= man_result_all_ones(8);
	wire_w_man_result_all_ones_range3473w(0) <= man_result_all_ones(9);
	wire_w_man_round_wi_range3474w(0) <= man_round_wi(10);
	wire_w_man_round_wi_range3477w(0) <= man_round_wi(11);
	wire_w_man_round_wi_range3480w(0) <= man_round_wi(12);
	wire_w_man_round_wi_range3483w(0) <= man_round_wi(13);
	wire_w_man_round_wi_range3486w(0) <= man_round_wi(14);
	wire_w_man_round_wi_range3489w(0) <= man_round_wi(15);
	wire_w_man_round_wi_range3492w(0) <= man_round_wi(16);
	wire_w_man_round_wi_range3495w(0) <= man_round_wi(17);
	wire_w_man_round_wi_range3498w(0) <= man_round_wi(18);
	wire_w_man_round_wi_range3501w(0) <= man_round_wi(19);
	wire_w_man_round_wi_range3447w(0) <= man_round_wi(1);
	wire_w_man_round_wi_range3504w(0) <= man_round_wi(20);
	wire_w_man_round_wi_range3507w(0) <= man_round_wi(21);
	wire_w_man_round_wi_range3510w(0) <= man_round_wi(22);
	wire_w_man_round_wi_range3513w(0) <= man_round_wi(23);
	wire_w_man_round_wi_range3516w(0) <= man_round_wi(24);
	wire_w_man_round_wi_range3519w(0) <= man_round_wi(25);
	wire_w_man_round_wi_range3522w(0) <= man_round_wi(26);
	wire_w_man_round_wi_range3525w(0) <= man_round_wi(27);
	wire_w_man_round_wi_range3528w(0) <= man_round_wi(28);
	wire_w_man_round_wi_range3531w(0) <= man_round_wi(29);
	wire_w_man_round_wi_range3450w(0) <= man_round_wi(2);
	wire_w_man_round_wi_range3534w(0) <= man_round_wi(30);
	wire_w_man_round_wi_range3537w(0) <= man_round_wi(31);
	wire_w_man_round_wi_range3540w(0) <= man_round_wi(32);
	wire_w_man_round_wi_range3543w(0) <= man_round_wi(33);
	wire_w_man_round_wi_range3546w(0) <= man_round_wi(34);
	wire_w_man_round_wi_range3549w(0) <= man_round_wi(35);
	wire_w_man_round_wi_range3552w(0) <= man_round_wi(36);
	wire_w_man_round_wi_range3555w(0) <= man_round_wi(37);
	wire_w_man_round_wi_range3558w(0) <= man_round_wi(38);
	wire_w_man_round_wi_range3561w(0) <= man_round_wi(39);
	wire_w_man_round_wi_range3453w(0) <= man_round_wi(3);
	wire_w_man_round_wi_range3564w(0) <= man_round_wi(40);
	wire_w_man_round_wi_range3567w(0) <= man_round_wi(41);
	wire_w_man_round_wi_range3570w(0) <= man_round_wi(42);
	wire_w_man_round_wi_range3573w(0) <= man_round_wi(43);
	wire_w_man_round_wi_range3576w(0) <= man_round_wi(44);
	wire_w_man_round_wi_range3579w(0) <= man_round_wi(45);
	wire_w_man_round_wi_range3582w(0) <= man_round_wi(46);
	wire_w_man_round_wi_range3585w(0) <= man_round_wi(47);
	wire_w_man_round_wi_range3588w(0) <= man_round_wi(48);
	wire_w_man_round_wi_range3591w(0) <= man_round_wi(49);
	wire_w_man_round_wi_range3456w(0) <= man_round_wi(4);
	wire_w_man_round_wi_range3594w(0) <= man_round_wi(50);
	wire_w_man_round_wi_range3597w(0) <= man_round_wi(51);
	wire_w_man_round_wi_range3459w(0) <= man_round_wi(5);
	wire_w_man_round_wi_range3462w(0) <= man_round_wi(6);
	wire_w_man_round_wi_range3465w(0) <= man_round_wi(7);
	wire_w_man_round_wi_range3468w(0) <= man_round_wi(8);
	wire_w_man_round_wi_range3471w(0) <= man_round_wi(9);
	wire_w_sticky_bits_range3395w(0) <= sticky_bits(0);
	wire_w_sticky_bits_range3399w(0) <= sticky_bits(1);
	wire_w_sticky_bits_range3402w(0) <= sticky_bits(2);
	wire_w_sticky_bits_range3405w(0) <= sticky_bits(3);
	wire_w_xf_pre_2_wo_range285w <= xf_pre_2_wo(59 DOWNTO 0);
	wire_w_xf_pre_wo_range279w <= xf_pre_wo(59 DOWNTO 0);
	man_prod :  ALTFP_EXa_altmult_opt_v4e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => tbl1_tbl2_prod_wo,
		datab => tbl3_taylor_prod_wo,
		result => wire_man_prod_result
	  );
	tbl1_tbl2_prod :  ALTFP_EXa_altmult_opt_45e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => table_one_out_pl,
		datab => table_two_out_pl,
		result => wire_tbl1_tbl2_prod_result
	  );
	wire_tbl3_taylor_prod_datab <= ( "1" & "000000000000000000000000000" & xf_pl(30 DOWNTO 0));
	tbl3_taylor_prod :  ALTFP_EXa_altmult_opt_95e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => table_three_out_pl,
		datab => wire_tbl3_taylor_prod_datab,
		result => wire_tbl3_taylor_prod_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes0 <= barrel_shifter_underflow_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes1 <= barrel_shifter_underflow_dffe2_23_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes2 <= barrel_shifter_underflow_dffe2_23_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes3 <= barrel_shifter_underflow_dffe2_23_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes4 <= barrel_shifter_underflow_dffe2_23_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes5 <= barrel_shifter_underflow_dffe2_23_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes6 <= barrel_shifter_underflow_dffe2_23_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes7 <= barrel_shifter_underflow_dffe2_23_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes8 <= barrel_shifter_underflow_dffe2_23_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes9 <= barrel_shifter_underflow_dffe2_23_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes10 <= barrel_shifter_underflow_dffe2_23_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes11 <= barrel_shifter_underflow_dffe2_23_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes12 <= barrel_shifter_underflow_dffe2_23_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes13 <= barrel_shifter_underflow_dffe2_23_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes14 <= barrel_shifter_underflow_dffe2_23_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes15 <= barrel_shifter_underflow_dffe2_23_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes16 <= barrel_shifter_underflow_dffe2_23_pipes15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes17 <= barrel_shifter_underflow_dffe2_23_pipes16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes18 <= barrel_shifter_underflow_dffe2_23_pipes17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes19 <= barrel_shifter_underflow_dffe2_23_pipes18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes20 <= barrel_shifter_underflow_dffe2_23_pipes19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes21 <= barrel_shifter_underflow_dffe2_23_pipes20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_23_pipes22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_23_pipes22 <= barrel_shifter_underflow_dffe2_23_pipes21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes0 <= distance_overflow_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes1 <= distance_overflow_dffe2_23_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes2 <= distance_overflow_dffe2_23_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes3 <= distance_overflow_dffe2_23_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes4 <= distance_overflow_dffe2_23_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes5 <= distance_overflow_dffe2_23_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes6 <= distance_overflow_dffe2_23_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes7 <= distance_overflow_dffe2_23_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes8 <= distance_overflow_dffe2_23_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes9 <= distance_overflow_dffe2_23_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes10 <= distance_overflow_dffe2_23_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes11 <= distance_overflow_dffe2_23_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes12 <= distance_overflow_dffe2_23_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes13 <= distance_overflow_dffe2_23_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes14 <= distance_overflow_dffe2_23_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes15 <= distance_overflow_dffe2_23_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes16 <= distance_overflow_dffe2_23_pipes15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes17 <= distance_overflow_dffe2_23_pipes16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes18 <= distance_overflow_dffe2_23_pipes17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes19 <= distance_overflow_dffe2_23_pipes18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes20 <= distance_overflow_dffe2_23_pipes19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes21 <= distance_overflow_dffe2_23_pipes20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_23_pipes22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_23_pipes22 <= distance_overflow_dffe2_23_pipes21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_0 <= wire_exp_value_b4_biasa_dataout;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_1 <= exp_value_b4_bias_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_10 <= exp_value_b4_bias_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_11 <= exp_value_b4_bias_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_12 <= exp_value_b4_bias_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_13 <= exp_value_b4_bias_dffe_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_14 <= exp_value_b4_bias_dffe_13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_15 <= exp_value_b4_bias_dffe_14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_16 <= exp_value_b4_bias_dffe_15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_17 <= exp_value_b4_bias_dffe_16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_18 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_18 <= exp_value_b4_bias_dffe_17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_2 <= exp_value_b4_bias_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_3 <= exp_value_b4_bias_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_4 <= exp_value_b4_bias_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_5 <= exp_value_b4_bias_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_6 <= exp_value_b4_bias_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_7 <= exp_value_b4_bias_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_8 <= exp_value_b4_bias_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_9 <= exp_value_b4_bias_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_dffe1 <= exp_value_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_0 <= extra_ln2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_1 <= extra_ln2_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_10 <= extra_ln2_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_11 <= extra_ln2_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	wire_extra_ln2_dffe_11_w_lg_q259w(0) <= NOT extra_ln2_dffe_11;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_2 <= extra_ln2_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_3 <= extra_ln2_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_4 <= extra_ln2_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_5 <= extra_ln2_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_6 <= extra_ln2_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_7 <= extra_ln2_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_8 <= extra_ln2_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_9 <= extra_ln2_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN fraction_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN fraction_dffe1 <= fraction_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes0 <= input_is_infinity_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes1 <= input_is_infinity_24_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes2 <= input_is_infinity_24_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes3 <= input_is_infinity_24_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes4 <= input_is_infinity_24_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes5 <= input_is_infinity_24_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes6 <= input_is_infinity_24_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes7 <= input_is_infinity_24_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes8 <= input_is_infinity_24_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes9 <= input_is_infinity_24_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes10 <= input_is_infinity_24_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes11 <= input_is_infinity_24_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes12 <= input_is_infinity_24_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes13 <= input_is_infinity_24_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes14 <= input_is_infinity_24_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes15 <= input_is_infinity_24_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes16 <= input_is_infinity_24_pipes15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes17 <= input_is_infinity_24_pipes16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes18 <= input_is_infinity_24_pipes17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes19 <= input_is_infinity_24_pipes18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes20 <= input_is_infinity_24_pipes19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes21 <= input_is_infinity_24_pipes20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes22 <= input_is_infinity_24_pipes21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_24_pipes23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_24_pipes23 <= input_is_infinity_24_pipes22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes0 <= input_is_nan_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes1 <= input_is_nan_24_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes2 <= input_is_nan_24_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes3 <= input_is_nan_24_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes4 <= input_is_nan_24_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes5 <= input_is_nan_24_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes6 <= input_is_nan_24_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes7 <= input_is_nan_24_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes8 <= input_is_nan_24_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes9 <= input_is_nan_24_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes10 <= input_is_nan_24_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes11 <= input_is_nan_24_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes12 <= input_is_nan_24_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes13 <= input_is_nan_24_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes14 <= input_is_nan_24_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes15 <= input_is_nan_24_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes16 <= input_is_nan_24_pipes15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes17 <= input_is_nan_24_pipes16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes18 <= input_is_nan_24_pipes17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes19 <= input_is_nan_24_pipes18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes20 <= input_is_nan_24_pipes19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes21 <= input_is_nan_24_pipes20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes22 <= input_is_nan_24_pipes21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_24_pipes23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_24_pipes23 <= input_is_nan_24_pipes22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes0 <= input_is_zero_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes1 <= input_is_zero_24_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes2 <= input_is_zero_24_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes3 <= input_is_zero_24_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes4 <= input_is_zero_24_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes5 <= input_is_zero_24_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes6 <= input_is_zero_24_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes7 <= input_is_zero_24_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes8 <= input_is_zero_24_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes9 <= input_is_zero_24_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes10 <= input_is_zero_24_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes11 <= input_is_zero_24_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes12 <= input_is_zero_24_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes13 <= input_is_zero_24_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes14 <= input_is_zero_24_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes15 <= input_is_zero_24_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes16 <= input_is_zero_24_pipes15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes17 <= input_is_zero_24_pipes16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes18 <= input_is_zero_24_pipes17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes19 <= input_is_zero_24_pipes18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes20 <= input_is_zero_24_pipes19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes21 <= input_is_zero_24_pipes20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes22 <= input_is_zero_24_pipes21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_24_pipes23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_24_pipes23 <= input_is_zero_24_pipes22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_overflow_dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_overflow_dffe15 <= man_overflow_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_round_dffe15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_round_dffe15 <= man_round_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_pipe_dffe16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_pipe_dffe16 <= result_pipe_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_up_dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_up_dffe15 <= round_up_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe0 <= sign_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe1 <= sign_dffe0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe2 <= sign_dffe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe3 <= sign_dffe2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe4 <= sign_dffe3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe5 <= sign_dffe4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe6 <= sign_dffe5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe7 <= sign_dffe6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe8 <= sign_dffe7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe9 <= sign_dffe8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe10 <= sign_dffe9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe11 <= sign_dffe10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe12 <= sign_dffe11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe13 <= sign_dffe12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe14 <= sign_dffe13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe15 <= sign_dffe14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe16 <= sign_dffe15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe17 <= sign_dffe16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe18 <= sign_dffe17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe19 <= sign_dffe18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe20 <= sign_dffe19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe21 <= sign_dffe20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe22 <= sign_dffe21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe23 <= sign_dffe22;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_dffe_w_lg_q3430w(0) <= sign_dffe23 AND wire_w_lg_distance_overflow3429w(0);
	wire_sign_dffe_w_lg_q3416w(0) <= NOT sign_dffe23;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN table_one_dffe12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN table_one_dffe12 <= table_one_out;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN table_three_dffe12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN table_three_dffe12 <= table_three_out;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN table_two_dffe12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN table_two_dffe12 <= table_two_out;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes0 <= tbl1_compare_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes1 <= tbl1_compare_dffe11_10_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes2 <= tbl1_compare_dffe11_10_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes3 <= tbl1_compare_dffe11_10_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes4 <= tbl1_compare_dffe11_10_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes5 <= tbl1_compare_dffe11_10_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes6 <= tbl1_compare_dffe11_10_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes7 <= tbl1_compare_dffe11_10_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes8 <= tbl1_compare_dffe11_10_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_10_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_10_pipes9 <= tbl1_compare_dffe11_10_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_0 <= x_fixed;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_1 <= x_fixed_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_2 <= x_fixed_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_3 <= x_fixed_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_4 <= x_fixed_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_5 <= x_fixed_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_6 <= x_fixed_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xf_pl_dffe12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xf_pl_dffe12 <= xf;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xf_pre_2_dffe10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xf_pre_2_dffe10 <= xf_pre_2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xf_pre_dffe9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xf_pre_dffe9 <= xf_pre_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xi_exp_value_dffe4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xi_exp_value_dffe4 <= xi_exp_value_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xi_ln2_prod_dffe7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xi_ln2_prod_dffe7 <= xi_ln2_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xi_prod_dffe3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xi_prod_dffe3 <= xi_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_minus_bias_dataa <= ( "0" & exp_w);
	wire_exp_minus_bias_datab <= ( "0" & exp_bias);
	exp_minus_bias :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => wire_exp_minus_bias_dataa,
		datab => wire_exp_minus_bias_datab,
		result => wire_exp_minus_bias_result
	  );
	wire_exp_value_add_bias_w_lg_w_result_range3427w3428w(0) <= NOT wire_exp_value_add_bias_w_result_range3427w(0);
	wire_exp_value_add_bias_dataa <= ( "0" & exp_value_b4_bias_dffe_18);
	wire_exp_value_add_bias_datab <= ( "0" & exp_bias(10 DOWNTO 1) & wire_extra_ln2_dffe_11_w_lg_q259w);
	wire_exp_value_add_bias_w_result_range3427w(0) <= wire_exp_value_add_bias_result(11);
	exp_value_add_bias :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_cin_to_bias_dataout,
		clken => clk_en,
		clock => clock,
		dataa => wire_exp_value_add_bias_dataa,
		datab => wire_exp_value_add_bias_datab,
		result => wire_exp_value_add_bias_result
	  );
	wire_exp_value_man_over_w_lg_w_lg_w_result_range3417w3418w3419w(0) <= wire_exp_value_man_over_w_lg_w_result_range3417w3418w(0) AND wire_sign_dffe_w_lg_q3416w(0);
	wire_exp_value_man_over_w_lg_w_result_range3417w3418w(0) <= NOT wire_exp_value_man_over_w_result_range3417w(0);
	wire_exp_value_man_over_w_lg_w_lg_w_lg_w_result_range3417w3418w3419w3420w(0) <= wire_exp_value_man_over_w_lg_w_lg_w_result_range3417w3418w3419w(0) OR sign_dffe23;
	wire_exp_value_man_over_datab <= ( "00000000000" & man_overflow_wo);
	wire_exp_value_man_over_w_result_range3417w(0) <= wire_exp_value_man_over_result(11);
	exp_value_man_over :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => wire_exp_value_add_bias_result,
		datab => wire_exp_value_man_over_datab,
		result => wire_exp_value_man_over_result
	  );
	wire_invert_exp_value_dataa <= (OTHERS => '0');
	wire_invert_exp_value_w_result_range232w <= wire_invert_exp_value_result(6 DOWNTO 0);
	invert_exp_value :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_invert_exp_value_dataa,
		datab => exp_value(10 DOWNTO 0),
		result => wire_invert_exp_value_result
	  );
	wire_man_round_datab <= ( "000000000000000000000000000000000000000000000000000" & round_up_wo);
	man_round :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 52
	  )
	  PORT MAP ( 
		dataa => man_round_wo,
		datab => wire_man_round_datab,
		result => wire_man_round_result
	  );
	wire_one_minus_xf_dataa <= ( "1" & "00000000000000000000000000000000000000000000000000000000000");
	one_minus_xf :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 60
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_one_minus_xf_dataa,
		datab => wire_extra_ln2_muxa_dataout,
		result => wire_one_minus_xf_result
	  );
	wire_x_fixed_minus_xiln2_datab <= ( "0" & xi_ln2_prod_wo(80 DOWNTO 12));
	x_fixed_minus_xiln2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 70
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => x_fixed_dffe_6,
		datab => wire_x_fixed_minus_xiln2_datab,
		result => wire_x_fixed_minus_xiln2_result
	  );
	wire_xf_minus_ln2_datab <= ( "00" & ln2_w(69 DOWNTO 12));
	xf_minus_ln2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 60
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => xf_pre(59 DOWNTO 0),
		datab => wire_xf_minus_ln2_datab,
		result => wire_xf_minus_ln2_result
	  );
	wire_xi_add_one_datab <= "00000000001";
	xi_add_one :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => xi_exp_value,
		datab => wire_xi_add_one_datab,
		result => wire_xi_add_one_result
	  );
	rbarrel_shift :  lpm_clshift
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_SHIFTTYPE => "LOGICAL",
		LPM_WIDTH => 70,
		LPM_WIDTHDIST => 7
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => barrel_shifter_data,
		direction => exp_value_wo(11),
		distance => barrel_shifter_distance,
		result => wire_rbarrel_shift_result
	  );
	distance_overflow_comp :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		agb => wire_distance_overflow_comp_agb,
		dataa => wire_exp_value_to_compare_muxa_dataout,
		datab => distance_overflow_val_w
	  );
	tbl1_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		ageb => wire_tbl1_compare_ageb,
		dataa => xf(57 DOWNTO 49),
		datab => addr_val_more_than_one
	  );
	underflow_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		agb => wire_underflow_compare_agb,
		dataa => wire_exp_value_to_compare_muxa_dataout,
		datab => underflow_compare_val_w
	  );
	xi_ln2_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 4,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 11,
		LPM_WIDTHB => 70,
		LPM_WIDTHP => 81,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_exp_value_to_ln2a_dataout,
		datab => ln2_w,
		result => wire_xi_ln2_prod_result
	  );
	xi_prod :  lpm_mult
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 15,
		LPM_WIDTHB => 12,
		LPM_WIDTHP => 27,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		dataa => x_fixed(69 DOWNTO 55),
		datab => one_over_ln2_w,
		result => wire_xi_prod_result
	  );
	loop2 : FOR i IN 0 TO 511 GENERATE
		loop3 : FOR j IN 0 TO 60 GENERATE
			wire_table_one_data_2d(i, j) <= table_one_data(i*61+j);
		END GENERATE loop3;
	END GENERATE loop2;
	table_one :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 512,
		LPM_WIDTH => 61,
		LPM_WIDTHS => 9
	  )
	  PORT MAP ( 
		data => wire_table_one_data_2d,
		result => wire_table_one_result,
		sel => xf(57 DOWNTO 49)
	  );
	loop4 : FOR i IN 0 TO 511 GENERATE
		loop5 : FOR j IN 0 TO 41 GENERATE
			wire_table_three_data_2d(i, j) <= table_three_data(i*42+j);
		END GENERATE loop5;
	END GENERATE loop4;
	table_three :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 512,
		LPM_WIDTH => 42,
		LPM_WIDTHS => 9
	  )
	  PORT MAP ( 
		data => wire_table_three_data_2d,
		result => wire_table_three_result,
		sel => xf(39 DOWNTO 31)
	  );
	loop6 : FOR i IN 0 TO 511 GENERATE
		loop7 : FOR j IN 0 TO 50 GENERATE
			wire_table_two_data_2d(i, j) <= table_two_data(i*51+j);
		END GENERATE loop7;
	END GENERATE loop6;
	table_two :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 512,
		LPM_WIDTH => 51,
		LPM_WIDTHS => 9
	  )
	  PORT MAP ( 
		data => wire_table_two_data_2d,
		result => wire_table_two_result,
		sel => xf(48 DOWNTO 40)
	  );
	wire_cin_to_bias_dataout <= shifted_value;
	wire_exp_result_mux_prea_dataout <= exp_one WHEN wire_w_lg_w3620w3621w(0) = '1'  ELSE exp_result_w;
	loop8 : FOR i IN 0 TO 10 GENERATE 
		wire_exp_result_mux_prea_w_lg_dataout3626w(i) <= wire_exp_result_mux_prea_dataout(i) AND wire_w_lg_w_lg_w_lg_underflow_w3623w3624w3625w(0);
	END GENERATE loop8;
	wire_exp_value_b4_biasa_dataout <= exp_invert WHEN sign_dffe3 = '1'  ELSE xi_exp_value;
	wire_exp_value_selecta_dataout <= wire_invert_exp_value_result(6 DOWNTO 0) WHEN exp_value_wo(11) = '1'  ELSE exp_value_wo(6 DOWNTO 0);
	wire_exp_value_to_compare_muxa_dataout <= wire_invert_exp_value_result WHEN exp_value_wo(11) = '1'  ELSE exp_value_wo(10 DOWNTO 0);
	wire_exp_value_to_ln2a_dataout <= wire_xi_add_one_result WHEN sign_dffe4 = '1'  ELSE xi_exp_value_wo;
	wire_extra_ln2_muxa_dataout <= wire_xf_minus_ln2_result WHEN extra_ln2_dffe_0 = '1'  ELSE xf_pre_wo(59 DOWNTO 0);
	wire_man_result_muxa_dataout <= ( nan_w & "000000000000000000000000000000000000000000000000000") WHEN wire_w_lg_w_lg_w_lg_w_lg_overflow_w3605w3606w3607w3608w(0) = '1'  ELSE wire_man_round_result;
	wire_xf_muxa_dataout <= wire_one_minus_xf_result WHEN sign_dffe12 = '1'  ELSE xf_pre_2_wo(59 DOWNTO 0);

 END RTL; --ALTFP_EXa_altfp_exp_iuc
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ALTFP_EXa IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END ALTFP_EXa;


ARCHITECTURE RTL OF altfp_exa IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (63 DOWNTO 0);



	COMPONENT ALTFP_EXa_altfp_exp_iuc
	PORT (
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(63 DOWNTO 0);

	ALTFP_EXa_altfp_exp_iuc_component : ALTFP_EXa_altfp_exp_iuc
	PORT MAP (
		aclr => aclr,
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_exp"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "25"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "11"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "52"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: data 0 0 64 0 INPUT NODEFVAL "data[63..0]"
-- Retrieval info: CONNECT: @data 0 0 64 0 data 0 0 64 0
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTFP_EXP.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTFP_EXP.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTFP_EXP.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTFP_EXP_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTFP_EXP.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTFP_EXP.cmp TRUE TRUE
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX NUMERIC "1"
-- Retrieval info: LIB_FILE: lpm
