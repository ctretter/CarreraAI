-------------------------------------------------------------------------------
-- Title      : Testbench for functions in global project package
-- Project    : Audio Signal Processing
-------------------------------------------------------------------------------
-- $Id: tbGlobal-e.vhd 3 2011-09-10 08:35:02Z mroland $
-------------------------------------------------------------------------------
-- Author     : Copyright 2003: Markus Pfaff
-- Standard   : Using VHDL'93
-- Simulation : Model Technology Modelsim
-- Synthesis  : Exemplar Leonardo
-------------------------------------------------------------------------------
-- Description:
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

use work.Global.all;

entity tbGlobal is

end entity tbGlobal;

