-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: tofixed.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.0.0 Build 211 04/27/2016 SJ Standard Edition
-- ************************************************************


--Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="FLOAT2FIXED" ROUNDING="TO_NEAREST" WIDTH_DATA=64 WIDTH_EXP_INPUT=11 WIDTH_EXP_OUTPUT=8 WIDTH_INT=12 WIDTH_MAN_INPUT=52 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=64 aclr clock dataa result
--VERSION_BEGIN 16.0 cbx_altbarrel_shift 2016:04:27:18:05:34:SJ cbx_altera_syncram_nd_impl 2016:04:27:18:05:34:SJ cbx_altfp_convert 2016:04:27:18:05:34:SJ cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_altsyncram 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_abs 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_decode 2016:04:27:18:05:34:SJ cbx_lpm_divide 2016:04:27:18:05:34:SJ cbx_lpm_mux 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_stratixiii 2016:04:27:18:05:34:SJ cbx_stratixv 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=2 SHIFTDIR="VARIABLE" SHIFTTYPE="LOGICAL" WIDTH=115 WIDTHDIST=7 aclr clk_en clock data direction distance result
--VERSION_BEGIN 16.0 cbx_altbarrel_shift 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END

--synthesis_resources = reg 235 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  tofixed_altbarrel_shift_v5h IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (114 DOWNTO 0);
		 direction	:	IN  STD_LOGIC := '0';
		 distance	:	IN  STD_LOGIC_VECTOR (6 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (114 DOWNTO 0)
	 ); 
 END tofixed_altbarrel_shift_v5h;

 ARCHITECTURE RTL OF tofixed_altbarrel_shift_v5h IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(114 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(114 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec5r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec6r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w527w528w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w523w524w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w548w549w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w544w545w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w570w571w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w566w567w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w592w593w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w588w589w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w614w615w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w610w611w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w633w634w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w629w630w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w654w655w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w650w651w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w519w520w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w540w541w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w562w563w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w584w585w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w606w607w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w625w626w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w646w647w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range515w527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range515w523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range536w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range536w544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range558w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range558w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range580w592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range580w588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range603w614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range603w610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range622w633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range622w629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range643w654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range643w650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range512w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range534w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range555w569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range577w591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range601w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range620w632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_dir_w_range640w653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range515w519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range536w540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range558w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range580w584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range603w606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range622w625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_sel_w_range643w646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range515w527w528w529w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range536w548w549w550w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range558w570w571w572w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range580w592w593w594w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range603w614w615w616w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range622w633w634w635w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range643w654w655w656w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w530w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w551w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w573w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w595w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w617w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w636w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w657w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (919 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (804 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w522w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w525w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w543w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w546w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w565w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w568w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w587w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w590w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w609w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w612w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w628w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w631w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w649w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w652w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_dir_w_range640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range510w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range533w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range553w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range575w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range597w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range619w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sbit_w_range638w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_sel_w_range643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_smux_w_range596w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_w_smux_w_range658w	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w527w528w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range515w527w(0) AND wire_altbarrel_shift2_w525w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w523w524w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range515w523w(0) AND wire_altbarrel_shift2_w522w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w548w549w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range536w548w(0) AND wire_altbarrel_shift2_w546w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w544w545w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range536w544w(0) AND wire_altbarrel_shift2_w543w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w570w571w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range558w570w(0) AND wire_altbarrel_shift2_w568w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w566w567w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range558w566w(0) AND wire_altbarrel_shift2_w565w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w592w593w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range580w592w(0) AND wire_altbarrel_shift2_w590w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w588w589w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range580w588w(0) AND wire_altbarrel_shift2_w587w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w614w615w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range603w614w(0) AND wire_altbarrel_shift2_w612w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w610w611w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range603w610w(0) AND wire_altbarrel_shift2_w609w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w633w634w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range622w633w(0) AND wire_altbarrel_shift2_w631w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w629w630w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range622w629w(0) AND wire_altbarrel_shift2_w628w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w654w655w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range643w654w(0) AND wire_altbarrel_shift2_w652w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w650w651w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range643w650w(0) AND wire_altbarrel_shift2_w649w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w519w520w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range515w519w(0) AND wire_altbarrel_shift2_w_sbit_w_range510w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w540w541w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range536w540w(0) AND wire_altbarrel_shift2_w_sbit_w_range533w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w562w563w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range558w562w(0) AND wire_altbarrel_shift2_w_sbit_w_range553w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w584w585w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range580w584w(0) AND wire_altbarrel_shift2_w_sbit_w_range575w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w606w607w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range603w606w(0) AND wire_altbarrel_shift2_w_sbit_w_range597w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w625w626w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range622w625w(0) AND wire_altbarrel_shift2_w_sbit_w_range619w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w646w647w(i) <= wire_altbarrel_shift2_w_lg_w_sel_w_range643w646w(0) AND wire_altbarrel_shift2_w_sbit_w_range638w(i);
	END GENERATE loop20;
	wire_altbarrel_shift2_w_lg_w_sel_w_range515w527w(0) <= wire_altbarrel_shift2_w_sel_w_range515w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range512w526w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range515w523w(0) <= wire_altbarrel_shift2_w_sel_w_range515w(0) AND wire_altbarrel_shift2_w_dir_w_range512w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range536w548w(0) <= wire_altbarrel_shift2_w_sel_w_range536w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range534w547w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range536w544w(0) <= wire_altbarrel_shift2_w_sel_w_range536w(0) AND wire_altbarrel_shift2_w_dir_w_range534w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range558w570w(0) <= wire_altbarrel_shift2_w_sel_w_range558w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range555w569w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range558w566w(0) <= wire_altbarrel_shift2_w_sel_w_range558w(0) AND wire_altbarrel_shift2_w_dir_w_range555w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range580w592w(0) <= wire_altbarrel_shift2_w_sel_w_range580w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range577w591w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range580w588w(0) <= wire_altbarrel_shift2_w_sel_w_range580w(0) AND wire_altbarrel_shift2_w_dir_w_range577w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range603w614w(0) <= wire_altbarrel_shift2_w_sel_w_range603w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range601w613w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range603w610w(0) <= wire_altbarrel_shift2_w_sel_w_range603w(0) AND wire_altbarrel_shift2_w_dir_w_range601w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range622w633w(0) <= wire_altbarrel_shift2_w_sel_w_range622w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range620w632w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range622w629w(0) <= wire_altbarrel_shift2_w_sel_w_range622w(0) AND wire_altbarrel_shift2_w_dir_w_range620w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range643w654w(0) <= wire_altbarrel_shift2_w_sel_w_range643w(0) AND wire_altbarrel_shift2_w_lg_w_dir_w_range640w653w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range643w650w(0) <= wire_altbarrel_shift2_w_sel_w_range643w(0) AND wire_altbarrel_shift2_w_dir_w_range640w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range512w526w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range512w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range534w547w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range534w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range555w569w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range555w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range577w591w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range577w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range601w613w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range601w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range620w632w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range620w(0);
	wire_altbarrel_shift2_w_lg_w_dir_w_range640w653w(0) <= NOT wire_altbarrel_shift2_w_dir_w_range640w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range515w519w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range515w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range536w540w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range536w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range558w562w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range558w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range580w584w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range580w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range603w606w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range603w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range622w625w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range622w(0);
	wire_altbarrel_shift2_w_lg_w_sel_w_range643w646w(0) <= NOT wire_altbarrel_shift2_w_sel_w_range643w(0);
	loop21 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range515w527w528w529w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w527w528w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w523w524w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range536w548w549w550w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w548w549w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w544w545w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range558w570w571w572w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w570w571w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w566w567w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range580w592w593w594w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w592w593w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w588w589w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range603w614w615w616w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w614w615w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w610w611w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range622w633w634w635w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w633w634w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w629w630w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range643w654w655w656w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w654w655w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w650w651w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w530w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range515w527w528w529w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range515w519w520w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w551w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range536w548w549w550w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range536w540w541w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w573w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range558w570w571w572w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range558w562w563w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w595w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range580w592w593w594w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range580w584w585w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w617w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range603w614w615w616w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range603w606w607w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w636w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range622w633w634w635w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range622w625w626w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 114 GENERATE 
		wire_altbarrel_shift2_w657w(i) <= wire_altbarrel_shift2_w_lg_w_lg_w_lg_w_sel_w_range643w654w655w656w(i) OR wire_altbarrel_shift2_w_lg_w_lg_w_sel_w_range643w646w647w(i);
	END GENERATE loop34;
	dir_w <= ( dir_pipe(1) & dir_w(5 DOWNTO 4) & dir_pipe(0) & dir_w(2 DOWNTO 0) & direction_w);
	direction_w <= direction;
	pad_w <= (OTHERS => '0');
	result <= sbit_w(919 DOWNTO 805);
	sbit_w <= ( sbit_piper2d & smux_w(689 DOWNTO 460) & sbit_piper1d & smux_w(344 DOWNTO 0) & data);
	sel_w <= ( sel_pipec6r1d & sel_pipec5r1d & sel_pipec4r1d & distance(3 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift2_w657w & wire_altbarrel_shift2_w636w & wire_altbarrel_shift2_w617w & wire_altbarrel_shift2_w595w & wire_altbarrel_shift2_w573w & wire_altbarrel_shift2_w551w & wire_altbarrel_shift2_w530w);
	wire_altbarrel_shift2_w522w <= ( pad_w(0) & sbit_w(114 DOWNTO 1));
	wire_altbarrel_shift2_w525w <= ( sbit_w(113 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift2_w543w <= ( pad_w(1 DOWNTO 0) & sbit_w(229 DOWNTO 117));
	wire_altbarrel_shift2_w546w <= ( sbit_w(227 DOWNTO 115) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift2_w565w <= ( pad_w(3 DOWNTO 0) & sbit_w(344 DOWNTO 234));
	wire_altbarrel_shift2_w568w <= ( sbit_w(340 DOWNTO 230) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift2_w587w <= ( pad_w(7 DOWNTO 0) & sbit_w(459 DOWNTO 353));
	wire_altbarrel_shift2_w590w <= ( sbit_w(451 DOWNTO 345) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift2_w609w <= ( pad_w(15 DOWNTO 0) & sbit_w(574 DOWNTO 476));
	wire_altbarrel_shift2_w612w <= ( sbit_w(558 DOWNTO 460) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift2_w628w <= ( pad_w(31 DOWNTO 0) & sbit_w(689 DOWNTO 607));
	wire_altbarrel_shift2_w631w <= ( sbit_w(657 DOWNTO 575) & pad_w(31 DOWNTO 0));
	wire_altbarrel_shift2_w649w <= ( pad_w(63 DOWNTO 0) & sbit_w(804 DOWNTO 754));
	wire_altbarrel_shift2_w652w <= ( sbit_w(740 DOWNTO 690) & pad_w(63 DOWNTO 0));
	wire_altbarrel_shift2_w_dir_w_range512w(0) <= dir_w(0);
	wire_altbarrel_shift2_w_dir_w_range534w(0) <= dir_w(1);
	wire_altbarrel_shift2_w_dir_w_range555w(0) <= dir_w(2);
	wire_altbarrel_shift2_w_dir_w_range577w(0) <= dir_w(3);
	wire_altbarrel_shift2_w_dir_w_range601w(0) <= dir_w(4);
	wire_altbarrel_shift2_w_dir_w_range620w(0) <= dir_w(5);
	wire_altbarrel_shift2_w_dir_w_range640w(0) <= dir_w(6);
	wire_altbarrel_shift2_w_sbit_w_range510w <= sbit_w(114 DOWNTO 0);
	wire_altbarrel_shift2_w_sbit_w_range533w <= sbit_w(229 DOWNTO 115);
	wire_altbarrel_shift2_w_sbit_w_range553w <= sbit_w(344 DOWNTO 230);
	wire_altbarrel_shift2_w_sbit_w_range575w <= sbit_w(459 DOWNTO 345);
	wire_altbarrel_shift2_w_sbit_w_range597w <= sbit_w(574 DOWNTO 460);
	wire_altbarrel_shift2_w_sbit_w_range619w <= sbit_w(689 DOWNTO 575);
	wire_altbarrel_shift2_w_sbit_w_range638w <= sbit_w(804 DOWNTO 690);
	wire_altbarrel_shift2_w_sel_w_range515w(0) <= sel_w(0);
	wire_altbarrel_shift2_w_sel_w_range536w(0) <= sel_w(1);
	wire_altbarrel_shift2_w_sel_w_range558w(0) <= sel_w(2);
	wire_altbarrel_shift2_w_sel_w_range580w(0) <= sel_w(3);
	wire_altbarrel_shift2_w_sel_w_range603w(0) <= sel_w(4);
	wire_altbarrel_shift2_w_sel_w_range622w(0) <= sel_w(5);
	wire_altbarrel_shift2_w_sel_w_range643w(0) <= sel_w(6);
	wire_altbarrel_shift2_w_smux_w_range596w <= smux_w(459 DOWNTO 345);
	wire_altbarrel_shift2_w_smux_w_range658w <= smux_w(804 DOWNTO 690);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(6) & dir_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift2_w_smux_w_range596w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift2_w_smux_w_range658w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec5r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec5r1d <= distance(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec6r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec6r1d <= distance(6);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --tofixed_altbarrel_shift_v5h

 LIBRARY lpm_ver;
 USE lpm_ver.all;

--synthesis_resources = lpm_add_sub 6 lpm_compare 4 reg 531 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  tofixed_altfp_convert_2gn IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END tofixed_altfp_convert_2gn;

 ARCHITECTURE RTL OF tofixed_altfp_convert_2gn IS

	 SIGNAL  wire_altbarrel_shift2_distance	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_barrel_direction_negative279w280w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift2_result	:	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL	 added_power2_reg	:	STD_LOGIC_VECTOR(6 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_direction_negative_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit3_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 border_lower_limit_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_border_lower_limit_reg4_w_lg_q489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_reg	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_equal_upper_limit_reg3_w_lg_q454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exceed_upper_limit_reg3_w_lg_q455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_or_reg4_w_lg_q220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 int_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_int_or_reg3_w_lg_q453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 integer_result_reg	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 integer_rounded_reg	:	STD_LOGIC_VECTOR(62 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_or_reg4_w_lg_q222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 mantissa_input_reg	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_exceeder_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 power2_value_reg	:	STD_LOGIC_VECTOR(6 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_input_reg3_w_lg_q456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sign_input_reg3_w_lg_q458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sign_input_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_adder_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_1_adder_datab	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_add_1_adder_result	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub3_w_lg_w_lg_cout465w466w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub3_w_lg_cout464w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub3_w_lg_cout465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub3_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub3_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub4_datab	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_barrel_direction_invert_dataa	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_barrel_direction_invert_result	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_lg_w_result_range257w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_lg_w_lg_w_result_range257w269w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_overflow	:	STD_LOGIC;
	 SIGNAL  wire_power2_value_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_power2_value_w_result_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_below_lower_limit1_aeb	:	STD_LOGIC;
	 SIGNAL  wire_below_lower_limit2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_exceed_upper_limit_aeb	:	STD_LOGIC;
	 SIGNAL  wire_exceed_upper_limit_agb	:	STD_LOGIC;
	 SIGNAL  wire_max_shift_compare_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_add_1_w441w442w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_barrel_direction_negative277w278w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_below_limit_exceeders495w496w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exceed_limit_exceeders506w507w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_lowest_integer_selector447w448w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w470w499w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w470w471w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w440w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_direction_negative279w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders494w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders505w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector446w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w498w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w469w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range228w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range232w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range235w237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range238w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range241w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range244w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range247w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range250w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range253w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_anding_range256w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range8w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range14w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range19w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range24w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range29w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range34w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range39w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range44w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range49w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range54w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_direction_negative277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_input_w501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_denormal_input_w490w491w492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_denormal_input_w490w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_infinity_input_w502w503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_denormal_input_w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinity_input_w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_oring_range260w262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_oring_range263w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_below_lower_limit3_oring_range265w266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range6w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range12w16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range17w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range22w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range27w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range32w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range37w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range42w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range47w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range52w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range108w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range105w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range102w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range99w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range96w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range93w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range90w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range87w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range84w86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range81w83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range135w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range78w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range75w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range72w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range69w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range66w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range62w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range132w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range129w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range126w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range123w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range120w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range117w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range114w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range111w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range187w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range184w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range181w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range178w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range175w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range172w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range169w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range166w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range163w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range160w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range214w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range157w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range154w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range151w153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range148w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range145w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range141w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range211w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range208w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range205w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range202w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range199w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range196w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range193w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range190w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range286w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range317w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range320w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range323w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range326w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range329w331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range332w334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range335w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range338w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range341w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range344w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range290w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range347w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range350w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range353w355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range356w358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range359w361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range362w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range365w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range368w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range371w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range374w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range293w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range377w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range380w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range383w385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range386w388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range389w391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range392w394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range395w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range398w400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range401w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range404w406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range296w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range407w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range410w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range413w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range416w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range419w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range422w424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range425w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range428w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range431w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range434w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range299w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range302w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range305w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range308w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range311w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range314w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_1_cout_w :	STD_LOGIC;
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  all_zeroes_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  barrel_direction_negative :	STD_LOGIC;
	 SIGNAL  barrel_mantissa_input :	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  barrel_zero_padding_w :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  below_limit_exceeders :	STD_LOGIC;
	 SIGNAL  below_limit_integer :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  below_lower_limit3_anding :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  below_lower_limit3_oring :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  below_lower_limit3_w :	STD_LOGIC;
	 SIGNAL  bias_value_less_1_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_res_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  denormal_input_w :	STD_LOGIC;
	 SIGNAL  equal_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exceed_limit_exceeders :	STD_LOGIC;
	 SIGNAL  exceed_limit_integer :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  exceed_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exp_and :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_and_w :	STD_LOGIC;
	 SIGNAL  exp_bus :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_or :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_or_w :	STD_LOGIC;
	 SIGNAL  exponent_input :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  implied_mantissa_input :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  infinity_input_w :	STD_LOGIC;
	 SIGNAL  infinity_value_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  int_or1_w :	STD_LOGIC;
	 SIGNAL  int_or2_w :	STD_LOGIC;
	 SIGNAL  integer_output :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  integer_post_round :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  integer_pre_round :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  integer_result :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  integer_rounded :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  integer_rounded_tmp :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  integer_tmp_output :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  inv_add_1_adder1_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  inv_add_1_adder2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  inv_integer :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  lbarrel_shift_result_w :	STD_LOGIC_VECTOR (114 DOWNTO 0);
	 SIGNAL  lbarrel_shift_w :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  lowest_integer_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_value :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  man_bus1 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_bus2 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_or1 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_or1_w :	STD_LOGIC;
	 SIGNAL  man_or2 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_or2_w :	STD_LOGIC;
	 SIGNAL  man_or_w :	STD_LOGIC;
	 SIGNAL  mantissa_input :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  max_shift_reg_w :	STD_LOGIC;
	 SIGNAL  max_shift_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  more_than_max_shift_w :	STD_LOGIC;
	 SIGNAL  nan_input_w :	STD_LOGIC;
	 SIGNAL  neg_infi_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  padded_exponent_input :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  pos_infi_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  power2_value_overflow_w :	STD_LOGIC;
	 SIGNAL  power2_value_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  shift_value_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  sign_input :	STD_LOGIC;
	 SIGNAL  sign_input_w :	STD_LOGIC;
	 SIGNAL  signed_integer :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  sticky_bus :	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  sticky_or :	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  unsigned_integer :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  upper_limit_w :	STD_LOGIC;
	 SIGNAL  zero_input_w :	STD_LOGIC;
	 SIGNAL  wire_w_below_lower_limit3_anding_range228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_anding_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_oring_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_oring_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_oring_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_below_lower_limit3_oring_range267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_inv_integer_range452w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  tofixed_altbarrel_shift_v5h
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(114 DOWNTO 0);
		direction	:	IN  STD_LOGIC := '0';
		distance	:	IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(114 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop35 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_w_lg_add_1_w441w442w(i) <= wire_w_lg_add_1_w441w(0) AND integer_pre_round(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_barrel_direction_negative277w278w(i) <= wire_w_lg_barrel_direction_negative277w(0) AND power2_value_reg(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 63 GENERATE 
		wire_w_lg_w_lg_below_limit_exceeders495w496w(i) <= wire_w_lg_below_limit_exceeders495w(0) AND integer_output(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 63 GENERATE 
		wire_w_lg_w_lg_exceed_limit_exceeders506w507w(i) <= wire_w_lg_exceed_limit_exceeders506w(0) AND below_limit_integer(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_w_lg_lowest_integer_selector447w448w(i) <= wire_w_lg_lowest_integer_selector447w(0) AND integer_rounded_tmp(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 63 GENERATE 
		wire_w_lg_w_lg_sign_input_w470w499w(i) <= wire_w_lg_sign_input_w470w(0) AND pos_infi_w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_w_lg_sign_input_w470w471w(i) <= wire_w_lg_sign_input_w470w(0) AND unsigned_integer(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_add_1_w440w(i) <= add_1_w AND integer_post_round(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_barrel_direction_negative279w(i) <= barrel_direction_negative AND wire_barrel_direction_invert_result(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 63 GENERATE 
		wire_w_lg_below_limit_exceeders494w(i) <= below_limit_exceeders AND all_zeroes_w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 63 GENERATE 
		wire_w_lg_exceed_limit_exceeders505w(i) <= exceed_limit_exceeders AND infinity_value_w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_lowest_integer_selector446w(i) <= lowest_integer_selector AND lowest_integer_value(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 63 GENERATE 
		wire_w_lg_sign_input_w498w(i) <= sign_input_w AND neg_infi_w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_sign_input_w469w(i) <= sign_input_w AND signed_integer(i);
	END GENERATE loop48;
	wire_w_lg_w_below_lower_limit3_anding_range228w231w(0) <= wire_w_below_lower_limit3_anding_range228w(0) AND wire_power2_value_w_result_range230w(0);
	wire_w_lg_w_below_lower_limit3_anding_range232w234w(0) <= wire_w_below_lower_limit3_anding_range232w(0) AND wire_power2_value_w_result_range233w(0);
	wire_w_lg_w_below_lower_limit3_anding_range235w237w(0) <= wire_w_below_lower_limit3_anding_range235w(0) AND wire_power2_value_w_result_range236w(0);
	wire_w_lg_w_below_lower_limit3_anding_range238w240w(0) <= wire_w_below_lower_limit3_anding_range238w(0) AND wire_power2_value_w_result_range239w(0);
	wire_w_lg_w_below_lower_limit3_anding_range241w243w(0) <= wire_w_below_lower_limit3_anding_range241w(0) AND wire_power2_value_w_result_range242w(0);
	wire_w_lg_w_below_lower_limit3_anding_range244w246w(0) <= wire_w_below_lower_limit3_anding_range244w(0) AND wire_power2_value_w_result_range245w(0);
	wire_w_lg_w_below_lower_limit3_anding_range247w249w(0) <= wire_w_below_lower_limit3_anding_range247w(0) AND wire_power2_value_w_result_range248w(0);
	wire_w_lg_w_below_lower_limit3_anding_range250w252w(0) <= wire_w_below_lower_limit3_anding_range250w(0) AND wire_power2_value_w_result_range251w(0);
	wire_w_lg_w_below_lower_limit3_anding_range253w255w(0) <= wire_w_below_lower_limit3_anding_range253w(0) AND wire_power2_value_w_result_range254w(0);
	wire_w_lg_w_below_lower_limit3_anding_range256w258w(0) <= wire_w_below_lower_limit3_anding_range256w(0) AND wire_power2_value_w_result_range257w(0);
	wire_w_lg_w_exp_and_range8w13w(0) <= wire_w_exp_and_range8w(0) AND wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_and_range14w18w(0) <= wire_w_exp_and_range14w(0) AND wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_and_range19w23w(0) <= wire_w_exp_and_range19w(0) AND wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_and_range24w28w(0) <= wire_w_exp_and_range24w(0) AND wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_and_range29w33w(0) <= wire_w_exp_and_range29w(0) AND wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_and_range34w38w(0) <= wire_w_exp_and_range34w(0) AND wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_and_range39w43w(0) <= wire_w_exp_and_range39w(0) AND wire_w_exp_bus_range40w(0);
	wire_w_lg_w_exp_and_range44w48w(0) <= wire_w_exp_and_range44w(0) AND wire_w_exp_bus_range45w(0);
	wire_w_lg_w_exp_and_range49w53w(0) <= wire_w_exp_and_range49w(0) AND wire_w_exp_bus_range50w(0);
	wire_w_lg_w_exp_and_range54w58w(0) <= wire_w_exp_and_range54w(0) AND wire_w_exp_bus_range55w(0);
	wire_w_lg_add_1_w441w(0) <= NOT add_1_w;
	wire_w_lg_barrel_direction_negative277w(0) <= NOT barrel_direction_negative;
	wire_w_lg_below_limit_exceeders495w(0) <= NOT below_limit_exceeders;
	wire_w_lg_exceed_limit_exceeders506w(0) <= NOT exceed_limit_exceeders;
	wire_w_lg_lowest_integer_selector447w(0) <= NOT lowest_integer_selector;
	wire_w_lg_nan_input_w501w(0) <= NOT nan_input_w;
	wire_w_lg_sign_input_w470w(0) <= NOT sign_input_w;
	wire_w_lg_w_lg_w_lg_denormal_input_w490w491w492w(0) <= wire_w_lg_w_lg_denormal_input_w490w491w(0) OR below_lower_limit3_reg4;
	wire_w_lg_w_lg_denormal_input_w490w491w(0) <= wire_w_lg_denormal_input_w490w(0) OR nan_input_w;
	wire_w_lg_w_lg_infinity_input_w502w503w(0) <= wire_w_lg_infinity_input_w502w(0) OR exceed_upper_limit_reg4;
	wire_w_lg_denormal_input_w490w(0) <= denormal_input_w OR zero_input_w;
	wire_w_lg_infinity_input_w502w(0) <= infinity_input_w OR max_shift_exceeder_reg;
	wire_w_lg_w_below_lower_limit3_oring_range260w262w(0) <= wire_w_below_lower_limit3_oring_range260w(0) OR wire_power2_value_w_result_range251w(0);
	wire_w_lg_w_below_lower_limit3_oring_range263w264w(0) <= wire_w_below_lower_limit3_oring_range263w(0) OR wire_power2_value_w_result_range254w(0);
	wire_w_lg_w_below_lower_limit3_oring_range265w266w(0) <= wire_w_below_lower_limit3_oring_range265w(0) OR wire_power2_value_w_result_range257w(0);
	wire_w_lg_w_exp_or_range6w11w(0) <= wire_w_exp_or_range6w(0) OR wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_or_range12w16w(0) <= wire_w_exp_or_range12w(0) OR wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_or_range17w21w(0) <= wire_w_exp_or_range17w(0) OR wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_or_range22w26w(0) <= wire_w_exp_or_range22w(0) OR wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_or_range27w31w(0) <= wire_w_exp_or_range27w(0) OR wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_or_range32w36w(0) <= wire_w_exp_or_range32w(0) OR wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_or_range37w41w(0) <= wire_w_exp_or_range37w(0) OR wire_w_exp_bus_range40w(0);
	wire_w_lg_w_exp_or_range42w46w(0) <= wire_w_exp_or_range42w(0) OR wire_w_exp_bus_range45w(0);
	wire_w_lg_w_exp_or_range47w51w(0) <= wire_w_exp_or_range47w(0) OR wire_w_exp_bus_range50w(0);
	wire_w_lg_w_exp_or_range52w56w(0) <= wire_w_exp_or_range52w(0) OR wire_w_exp_bus_range55w(0);
	wire_w_lg_w_man_or1_range108w110w(0) <= wire_w_man_or1_range108w(0) OR wire_w_man_bus1_range109w(0);
	wire_w_lg_w_man_or1_range105w107w(0) <= wire_w_man_or1_range105w(0) OR wire_w_man_bus1_range106w(0);
	wire_w_lg_w_man_or1_range102w104w(0) <= wire_w_man_or1_range102w(0) OR wire_w_man_bus1_range103w(0);
	wire_w_lg_w_man_or1_range99w101w(0) <= wire_w_man_or1_range99w(0) OR wire_w_man_bus1_range100w(0);
	wire_w_lg_w_man_or1_range96w98w(0) <= wire_w_man_or1_range96w(0) OR wire_w_man_bus1_range97w(0);
	wire_w_lg_w_man_or1_range93w95w(0) <= wire_w_man_or1_range93w(0) OR wire_w_man_bus1_range94w(0);
	wire_w_lg_w_man_or1_range90w92w(0) <= wire_w_man_or1_range90w(0) OR wire_w_man_bus1_range91w(0);
	wire_w_lg_w_man_or1_range87w89w(0) <= wire_w_man_or1_range87w(0) OR wire_w_man_bus1_range88w(0);
	wire_w_lg_w_man_or1_range84w86w(0) <= wire_w_man_or1_range84w(0) OR wire_w_man_bus1_range85w(0);
	wire_w_lg_w_man_or1_range81w83w(0) <= wire_w_man_or1_range81w(0) OR wire_w_man_bus1_range82w(0);
	wire_w_lg_w_man_or1_range135w137w(0) <= wire_w_man_or1_range135w(0) OR wire_w_man_bus1_range136w(0);
	wire_w_lg_w_man_or1_range78w80w(0) <= wire_w_man_or1_range78w(0) OR wire_w_man_bus1_range79w(0);
	wire_w_lg_w_man_or1_range75w77w(0) <= wire_w_man_or1_range75w(0) OR wire_w_man_bus1_range76w(0);
	wire_w_lg_w_man_or1_range72w74w(0) <= wire_w_man_or1_range72w(0) OR wire_w_man_bus1_range73w(0);
	wire_w_lg_w_man_or1_range69w71w(0) <= wire_w_man_or1_range69w(0) OR wire_w_man_bus1_range70w(0);
	wire_w_lg_w_man_or1_range66w68w(0) <= wire_w_man_or1_range66w(0) OR wire_w_man_bus1_range67w(0);
	wire_w_lg_w_man_or1_range62w65w(0) <= wire_w_man_or1_range62w(0) OR wire_w_man_bus1_range64w(0);
	wire_w_lg_w_man_or1_range132w134w(0) <= wire_w_man_or1_range132w(0) OR wire_w_man_bus1_range133w(0);
	wire_w_lg_w_man_or1_range129w131w(0) <= wire_w_man_or1_range129w(0) OR wire_w_man_bus1_range130w(0);
	wire_w_lg_w_man_or1_range126w128w(0) <= wire_w_man_or1_range126w(0) OR wire_w_man_bus1_range127w(0);
	wire_w_lg_w_man_or1_range123w125w(0) <= wire_w_man_or1_range123w(0) OR wire_w_man_bus1_range124w(0);
	wire_w_lg_w_man_or1_range120w122w(0) <= wire_w_man_or1_range120w(0) OR wire_w_man_bus1_range121w(0);
	wire_w_lg_w_man_or1_range117w119w(0) <= wire_w_man_or1_range117w(0) OR wire_w_man_bus1_range118w(0);
	wire_w_lg_w_man_or1_range114w116w(0) <= wire_w_man_or1_range114w(0) OR wire_w_man_bus1_range115w(0);
	wire_w_lg_w_man_or1_range111w113w(0) <= wire_w_man_or1_range111w(0) OR wire_w_man_bus1_range112w(0);
	wire_w_lg_w_man_or2_range187w189w(0) <= wire_w_man_or2_range187w(0) OR wire_w_man_bus2_range188w(0);
	wire_w_lg_w_man_or2_range184w186w(0) <= wire_w_man_or2_range184w(0) OR wire_w_man_bus2_range185w(0);
	wire_w_lg_w_man_or2_range181w183w(0) <= wire_w_man_or2_range181w(0) OR wire_w_man_bus2_range182w(0);
	wire_w_lg_w_man_or2_range178w180w(0) <= wire_w_man_or2_range178w(0) OR wire_w_man_bus2_range179w(0);
	wire_w_lg_w_man_or2_range175w177w(0) <= wire_w_man_or2_range175w(0) OR wire_w_man_bus2_range176w(0);
	wire_w_lg_w_man_or2_range172w174w(0) <= wire_w_man_or2_range172w(0) OR wire_w_man_bus2_range173w(0);
	wire_w_lg_w_man_or2_range169w171w(0) <= wire_w_man_or2_range169w(0) OR wire_w_man_bus2_range170w(0);
	wire_w_lg_w_man_or2_range166w168w(0) <= wire_w_man_or2_range166w(0) OR wire_w_man_bus2_range167w(0);
	wire_w_lg_w_man_or2_range163w165w(0) <= wire_w_man_or2_range163w(0) OR wire_w_man_bus2_range164w(0);
	wire_w_lg_w_man_or2_range160w162w(0) <= wire_w_man_or2_range160w(0) OR wire_w_man_bus2_range161w(0);
	wire_w_lg_w_man_or2_range214w216w(0) <= wire_w_man_or2_range214w(0) OR wire_w_man_bus2_range215w(0);
	wire_w_lg_w_man_or2_range157w159w(0) <= wire_w_man_or2_range157w(0) OR wire_w_man_bus2_range158w(0);
	wire_w_lg_w_man_or2_range154w156w(0) <= wire_w_man_or2_range154w(0) OR wire_w_man_bus2_range155w(0);
	wire_w_lg_w_man_or2_range151w153w(0) <= wire_w_man_or2_range151w(0) OR wire_w_man_bus2_range152w(0);
	wire_w_lg_w_man_or2_range148w150w(0) <= wire_w_man_or2_range148w(0) OR wire_w_man_bus2_range149w(0);
	wire_w_lg_w_man_or2_range145w147w(0) <= wire_w_man_or2_range145w(0) OR wire_w_man_bus2_range146w(0);
	wire_w_lg_w_man_or2_range141w144w(0) <= wire_w_man_or2_range141w(0) OR wire_w_man_bus2_range143w(0);
	wire_w_lg_w_man_or2_range211w213w(0) <= wire_w_man_or2_range211w(0) OR wire_w_man_bus2_range212w(0);
	wire_w_lg_w_man_or2_range208w210w(0) <= wire_w_man_or2_range208w(0) OR wire_w_man_bus2_range209w(0);
	wire_w_lg_w_man_or2_range205w207w(0) <= wire_w_man_or2_range205w(0) OR wire_w_man_bus2_range206w(0);
	wire_w_lg_w_man_or2_range202w204w(0) <= wire_w_man_or2_range202w(0) OR wire_w_man_bus2_range203w(0);
	wire_w_lg_w_man_or2_range199w201w(0) <= wire_w_man_or2_range199w(0) OR wire_w_man_bus2_range200w(0);
	wire_w_lg_w_man_or2_range196w198w(0) <= wire_w_man_or2_range196w(0) OR wire_w_man_bus2_range197w(0);
	wire_w_lg_w_man_or2_range193w195w(0) <= wire_w_man_or2_range193w(0) OR wire_w_man_bus2_range194w(0);
	wire_w_lg_w_man_or2_range190w192w(0) <= wire_w_man_or2_range190w(0) OR wire_w_man_bus2_range191w(0);
	wire_w_lg_w_sticky_or_range286w289w(0) <= wire_w_sticky_or_range286w(0) OR wire_w_sticky_bus_range288w(0);
	wire_w_lg_w_sticky_or_range317w319w(0) <= wire_w_sticky_or_range317w(0) OR wire_w_sticky_bus_range318w(0);
	wire_w_lg_w_sticky_or_range320w322w(0) <= wire_w_sticky_or_range320w(0) OR wire_w_sticky_bus_range321w(0);
	wire_w_lg_w_sticky_or_range323w325w(0) <= wire_w_sticky_or_range323w(0) OR wire_w_sticky_bus_range324w(0);
	wire_w_lg_w_sticky_or_range326w328w(0) <= wire_w_sticky_or_range326w(0) OR wire_w_sticky_bus_range327w(0);
	wire_w_lg_w_sticky_or_range329w331w(0) <= wire_w_sticky_or_range329w(0) OR wire_w_sticky_bus_range330w(0);
	wire_w_lg_w_sticky_or_range332w334w(0) <= wire_w_sticky_or_range332w(0) OR wire_w_sticky_bus_range333w(0);
	wire_w_lg_w_sticky_or_range335w337w(0) <= wire_w_sticky_or_range335w(0) OR wire_w_sticky_bus_range336w(0);
	wire_w_lg_w_sticky_or_range338w340w(0) <= wire_w_sticky_or_range338w(0) OR wire_w_sticky_bus_range339w(0);
	wire_w_lg_w_sticky_or_range341w343w(0) <= wire_w_sticky_or_range341w(0) OR wire_w_sticky_bus_range342w(0);
	wire_w_lg_w_sticky_or_range344w346w(0) <= wire_w_sticky_or_range344w(0) OR wire_w_sticky_bus_range345w(0);
	wire_w_lg_w_sticky_or_range290w292w(0) <= wire_w_sticky_or_range290w(0) OR wire_w_sticky_bus_range291w(0);
	wire_w_lg_w_sticky_or_range347w349w(0) <= wire_w_sticky_or_range347w(0) OR wire_w_sticky_bus_range348w(0);
	wire_w_lg_w_sticky_or_range350w352w(0) <= wire_w_sticky_or_range350w(0) OR wire_w_sticky_bus_range351w(0);
	wire_w_lg_w_sticky_or_range353w355w(0) <= wire_w_sticky_or_range353w(0) OR wire_w_sticky_bus_range354w(0);
	wire_w_lg_w_sticky_or_range356w358w(0) <= wire_w_sticky_or_range356w(0) OR wire_w_sticky_bus_range357w(0);
	wire_w_lg_w_sticky_or_range359w361w(0) <= wire_w_sticky_or_range359w(0) OR wire_w_sticky_bus_range360w(0);
	wire_w_lg_w_sticky_or_range362w364w(0) <= wire_w_sticky_or_range362w(0) OR wire_w_sticky_bus_range363w(0);
	wire_w_lg_w_sticky_or_range365w367w(0) <= wire_w_sticky_or_range365w(0) OR wire_w_sticky_bus_range366w(0);
	wire_w_lg_w_sticky_or_range368w370w(0) <= wire_w_sticky_or_range368w(0) OR wire_w_sticky_bus_range369w(0);
	wire_w_lg_w_sticky_or_range371w373w(0) <= wire_w_sticky_or_range371w(0) OR wire_w_sticky_bus_range372w(0);
	wire_w_lg_w_sticky_or_range374w376w(0) <= wire_w_sticky_or_range374w(0) OR wire_w_sticky_bus_range375w(0);
	wire_w_lg_w_sticky_or_range293w295w(0) <= wire_w_sticky_or_range293w(0) OR wire_w_sticky_bus_range294w(0);
	wire_w_lg_w_sticky_or_range377w379w(0) <= wire_w_sticky_or_range377w(0) OR wire_w_sticky_bus_range378w(0);
	wire_w_lg_w_sticky_or_range380w382w(0) <= wire_w_sticky_or_range380w(0) OR wire_w_sticky_bus_range381w(0);
	wire_w_lg_w_sticky_or_range383w385w(0) <= wire_w_sticky_or_range383w(0) OR wire_w_sticky_bus_range384w(0);
	wire_w_lg_w_sticky_or_range386w388w(0) <= wire_w_sticky_or_range386w(0) OR wire_w_sticky_bus_range387w(0);
	wire_w_lg_w_sticky_or_range389w391w(0) <= wire_w_sticky_or_range389w(0) OR wire_w_sticky_bus_range390w(0);
	wire_w_lg_w_sticky_or_range392w394w(0) <= wire_w_sticky_or_range392w(0) OR wire_w_sticky_bus_range393w(0);
	wire_w_lg_w_sticky_or_range395w397w(0) <= wire_w_sticky_or_range395w(0) OR wire_w_sticky_bus_range396w(0);
	wire_w_lg_w_sticky_or_range398w400w(0) <= wire_w_sticky_or_range398w(0) OR wire_w_sticky_bus_range399w(0);
	wire_w_lg_w_sticky_or_range401w403w(0) <= wire_w_sticky_or_range401w(0) OR wire_w_sticky_bus_range402w(0);
	wire_w_lg_w_sticky_or_range404w406w(0) <= wire_w_sticky_or_range404w(0) OR wire_w_sticky_bus_range405w(0);
	wire_w_lg_w_sticky_or_range296w298w(0) <= wire_w_sticky_or_range296w(0) OR wire_w_sticky_bus_range297w(0);
	wire_w_lg_w_sticky_or_range407w409w(0) <= wire_w_sticky_or_range407w(0) OR wire_w_sticky_bus_range408w(0);
	wire_w_lg_w_sticky_or_range410w412w(0) <= wire_w_sticky_or_range410w(0) OR wire_w_sticky_bus_range411w(0);
	wire_w_lg_w_sticky_or_range413w415w(0) <= wire_w_sticky_or_range413w(0) OR wire_w_sticky_bus_range414w(0);
	wire_w_lg_w_sticky_or_range416w418w(0) <= wire_w_sticky_or_range416w(0) OR wire_w_sticky_bus_range417w(0);
	wire_w_lg_w_sticky_or_range419w421w(0) <= wire_w_sticky_or_range419w(0) OR wire_w_sticky_bus_range420w(0);
	wire_w_lg_w_sticky_or_range422w424w(0) <= wire_w_sticky_or_range422w(0) OR wire_w_sticky_bus_range423w(0);
	wire_w_lg_w_sticky_or_range425w427w(0) <= wire_w_sticky_or_range425w(0) OR wire_w_sticky_bus_range426w(0);
	wire_w_lg_w_sticky_or_range428w430w(0) <= wire_w_sticky_or_range428w(0) OR wire_w_sticky_bus_range429w(0);
	wire_w_lg_w_sticky_or_range431w433w(0) <= wire_w_sticky_or_range431w(0) OR wire_w_sticky_bus_range432w(0);
	wire_w_lg_w_sticky_or_range434w436w(0) <= wire_w_sticky_or_range434w(0) OR wire_w_sticky_bus_range435w(0);
	wire_w_lg_w_sticky_or_range299w301w(0) <= wire_w_sticky_or_range299w(0) OR wire_w_sticky_bus_range300w(0);
	wire_w_lg_w_sticky_or_range302w304w(0) <= wire_w_sticky_or_range302w(0) OR wire_w_sticky_bus_range303w(0);
	wire_w_lg_w_sticky_or_range305w307w(0) <= wire_w_sticky_or_range305w(0) OR wire_w_sticky_bus_range306w(0);
	wire_w_lg_w_sticky_or_range308w310w(0) <= wire_w_sticky_or_range308w(0) OR wire_w_sticky_bus_range309w(0);
	wire_w_lg_w_sticky_or_range311w313w(0) <= wire_w_sticky_or_range311w(0) OR wire_w_sticky_bus_range312w(0);
	wire_w_lg_w_sticky_or_range314w316w(0) <= wire_w_sticky_or_range314w(0) OR wire_w_sticky_bus_range315w(0);
	add_1_cout_w <= ((wire_add_1_adder_cout AND add_1_w) AND wire_sign_input_reg3_w_lg_q458w(0));
	add_1_w <= (round_bit_w AND (guard_bit_w OR sticky_bit_w));
	all_zeroes_w <= ( "0" & "000000000000000000000000000000000000000000000000000000000000000");
	barrel_direction_negative <= barrel_direction_negative_reg;
	barrel_mantissa_input <= ( barrel_zero_padding_w & implied_mantissa_input);
	barrel_zero_padding_w <= (OTHERS => '0');
	below_limit_exceeders <= (wire_w_lg_w_lg_w_lg_denormal_input_w490w491w492w(0) AND wire_border_lower_limit_reg4_w_lg_q489w(0));
	below_limit_integer <= (wire_w_lg_w_lg_below_limit_exceeders495w496w OR wire_w_lg_below_limit_exceeders494w);
	below_lower_limit3_anding <= ( wire_w_lg_w_below_lower_limit3_anding_range256w258w & wire_w_lg_w_below_lower_limit3_anding_range253w255w & wire_w_lg_w_below_lower_limit3_anding_range250w252w & wire_w_lg_w_below_lower_limit3_anding_range247w249w & wire_w_lg_w_below_lower_limit3_anding_range244w246w & wire_w_lg_w_below_lower_limit3_anding_range241w243w & wire_w_lg_w_below_lower_limit3_anding_range238w240w & wire_w_lg_w_below_lower_limit3_anding_range235w237w & wire_w_lg_w_below_lower_limit3_anding_range232w234w & wire_w_lg_w_below_lower_limit3_anding_range228w231w & wire_power2_value_result(0));
	below_lower_limit3_oring <= ( wire_w_lg_w_below_lower_limit3_oring_range265w266w & wire_w_lg_w_below_lower_limit3_oring_range263w264w & wire_w_lg_w_below_lower_limit3_oring_range260w262w & wire_power2_value_result(7));
	below_lower_limit3_w <= (wire_power2_value_w_lg_w_lg_w_result_range257w269w270w(0) AND (NOT below_lower_limit3_anding(10)));
	bias_value_less_1_w <= "01111111110";
	clk_en <= '1';
	const_bias_value_add_width_res_w <= "10000001010";
	denormal_input_w <= (wire_exp_or_reg4_w_lg_q220w(0) AND man_or_reg4);
	equal_upper_limit_w <= wire_exceed_upper_limit_aeb;
	exceed_limit_exceeders <= (wire_w_lg_w_lg_infinity_input_w502w503w(0) AND wire_w_lg_nan_input_w501w(0));
	exceed_limit_integer <= (wire_w_lg_w_lg_exceed_limit_exceeders506w507w OR wire_w_lg_exceed_limit_exceeders505w);
	exceed_upper_limit_w <= wire_exceed_upper_limit_agb;
	exp_and <= ( wire_w_lg_w_exp_and_range54w58w & wire_w_lg_w_exp_and_range49w53w & wire_w_lg_w_exp_and_range44w48w & wire_w_lg_w_exp_and_range39w43w & wire_w_lg_w_exp_and_range34w38w & wire_w_lg_w_exp_and_range29w33w & wire_w_lg_w_exp_and_range24w28w & wire_w_lg_w_exp_and_range19w23w & wire_w_lg_w_exp_and_range14w18w & wire_w_lg_w_exp_and_range8w13w & exp_bus(0));
	exp_and_w <= exp_and(10);
	exp_bus <= exponent_input;
	exp_or <= ( wire_w_lg_w_exp_or_range52w56w & wire_w_lg_w_exp_or_range47w51w & wire_w_lg_w_exp_or_range42w46w & wire_w_lg_w_exp_or_range37w41w & wire_w_lg_w_exp_or_range32w36w & wire_w_lg_w_exp_or_range27w31w & wire_w_lg_w_exp_or_range22w26w & wire_w_lg_w_exp_or_range17w21w & wire_w_lg_w_exp_or_range12w16w & wire_w_lg_w_exp_or_range6w11w & exp_bus(0));
	exp_or_w <= exp_or(10);
	exponent_input <= dataa_reg(62 DOWNTO 52);
	guard_bit_w <= wire_altbarrel_shift2_result(52);
	implied_mantissa_input <= ( "1" & mantissa_input_reg);
	infinity_input_w <= (exp_and_reg4 AND wire_man_or_reg4_w_lg_q222w(0));
	infinity_value_w <= (wire_w_lg_w_lg_sign_input_w470w499w OR wire_w_lg_sign_input_w498w);
	int_or1_w <= man_or2(0);
	int_or2_w <= man_or1(0);
	integer_output <= ( sign_input_w & integer_tmp_output);
	integer_post_round <= wire_add_1_adder_result;
	integer_pre_round <= lbarrel_shift_w;
	integer_result <= exceed_limit_integer;
	integer_rounded <= (wire_w_lg_w_lg_lowest_integer_selector447w448w OR wire_w_lg_lowest_integer_selector446w);
	integer_rounded_tmp <= (wire_w_lg_w_lg_add_1_w441w442w OR wire_w_lg_add_1_w440w);
	integer_tmp_output <= (wire_w_lg_w_lg_sign_input_w470w471w OR wire_w_lg_sign_input_w469w);
	inv_add_1_adder1_w <= wire_add_sub3_result;
	inv_add_1_adder2_w <= (wire_add_sub3_w_lg_w_lg_cout465w466w OR wire_add_sub3_w_lg_cout464w);
	inv_integer <= (NOT integer_rounded_reg);
	lbarrel_shift_result_w <= wire_altbarrel_shift2_result;
	lbarrel_shift_w <= lbarrel_shift_result_w(114 DOWNTO 52);
	lowest_integer_selector <= '0';
	lowest_integer_value <= ( barrel_zero_padding_w & "1");
	man_bus1 <= mantissa_input(25 DOWNTO 0);
	man_bus2 <= mantissa_input(51 DOWNTO 26);
	man_or1 <= ( man_bus1(25) & wire_w_lg_w_man_or1_range62w65w & wire_w_lg_w_man_or1_range66w68w & wire_w_lg_w_man_or1_range69w71w & wire_w_lg_w_man_or1_range72w74w & wire_w_lg_w_man_or1_range75w77w & wire_w_lg_w_man_or1_range78w80w & wire_w_lg_w_man_or1_range81w83w & wire_w_lg_w_man_or1_range84w86w & wire_w_lg_w_man_or1_range87w89w & wire_w_lg_w_man_or1_range90w92w & wire_w_lg_w_man_or1_range93w95w & wire_w_lg_w_man_or1_range96w98w & wire_w_lg_w_man_or1_range99w101w & wire_w_lg_w_man_or1_range102w104w & wire_w_lg_w_man_or1_range105w107w & wire_w_lg_w_man_or1_range108w110w & wire_w_lg_w_man_or1_range111w113w & wire_w_lg_w_man_or1_range114w116w & wire_w_lg_w_man_or1_range117w119w & wire_w_lg_w_man_or1_range120w122w & wire_w_lg_w_man_or1_range123w125w & wire_w_lg_w_man_or1_range126w128w & wire_w_lg_w_man_or1_range129w131w & wire_w_lg_w_man_or1_range132w134w & wire_w_lg_w_man_or1_range135w137w);
	man_or1_w <= man_or1(0);
	man_or2 <= ( man_bus2(25) & wire_w_lg_w_man_or2_range141w144w & wire_w_lg_w_man_or2_range145w147w & wire_w_lg_w_man_or2_range148w150w & wire_w_lg_w_man_or2_range151w153w & wire_w_lg_w_man_or2_range154w156w & wire_w_lg_w_man_or2_range157w159w & wire_w_lg_w_man_or2_range160w162w & wire_w_lg_w_man_or2_range163w165w & wire_w_lg_w_man_or2_range166w168w & wire_w_lg_w_man_or2_range169w171w & wire_w_lg_w_man_or2_range172w174w & wire_w_lg_w_man_or2_range175w177w & wire_w_lg_w_man_or2_range178w180w & wire_w_lg_w_man_or2_range181w183w & wire_w_lg_w_man_or2_range184w186w & wire_w_lg_w_man_or2_range187w189w & wire_w_lg_w_man_or2_range190w192w & wire_w_lg_w_man_or2_range193w195w & wire_w_lg_w_man_or2_range196w198w & wire_w_lg_w_man_or2_range199w201w & wire_w_lg_w_man_or2_range202w204w & wire_w_lg_w_man_or2_range205w207w & wire_w_lg_w_man_or2_range208w210w & wire_w_lg_w_man_or2_range211w213w & wire_w_lg_w_man_or2_range214w216w);
	man_or2_w <= man_or2(0);
	man_or_w <= (man_or1_reg1 OR man_or2_reg1);
	mantissa_input <= dataa_reg(51 DOWNTO 0);
	max_shift_reg_w <= max_shift_reg;
	max_shift_w <= "0001010";
	more_than_max_shift_w <= (max_shift_reg_w AND add_1_cout_w);
	nan_input_w <= (exp_and_reg4 AND man_or_reg4);
	neg_infi_w <= ( "1" & "000000000000000000000000000000000000000000000000000000000000000");
	padded_exponent_input <= exponent_input;
	pos_infi_w <= ( "0" & "111111111111111111111111111111111111111111111111111111111111111");
	power2_value_overflow_w <= wire_power2_value_overflow;
	power2_value_w <= wire_power2_value_result(6 DOWNTO 0);
	result <= result_w;
	result_w <= integer_result_reg;
	round_bit_w <= wire_altbarrel_shift2_result(51);
	shift_value_w <= "01111001011";
	sign_input <= dataa_reg(63);
	sign_input_w <= sign_input_reg4;
	signed_integer <= ( inv_add_1_adder2_w & inv_add_1_adder1_w);
	sticky_bit_w <= sticky_or(50);
	sticky_bus <= wire_altbarrel_shift2_result(50 DOWNTO 0);
	sticky_or <= ( wire_w_lg_w_sticky_or_range434w436w & wire_w_lg_w_sticky_or_range431w433w & wire_w_lg_w_sticky_or_range428w430w & wire_w_lg_w_sticky_or_range425w427w & wire_w_lg_w_sticky_or_range422w424w & wire_w_lg_w_sticky_or_range419w421w & wire_w_lg_w_sticky_or_range416w418w & wire_w_lg_w_sticky_or_range413w415w & wire_w_lg_w_sticky_or_range410w412w & wire_w_lg_w_sticky_or_range407w409w & wire_w_lg_w_sticky_or_range404w406w & wire_w_lg_w_sticky_or_range401w403w & wire_w_lg_w_sticky_or_range398w400w & wire_w_lg_w_sticky_or_range395w397w & wire_w_lg_w_sticky_or_range392w394w & wire_w_lg_w_sticky_or_range389w391w & wire_w_lg_w_sticky_or_range386w388w & wire_w_lg_w_sticky_or_range383w385w & wire_w_lg_w_sticky_or_range380w382w & wire_w_lg_w_sticky_or_range377w379w & wire_w_lg_w_sticky_or_range374w376w & wire_w_lg_w_sticky_or_range371w373w & wire_w_lg_w_sticky_or_range368w370w & wire_w_lg_w_sticky_or_range365w367w & wire_w_lg_w_sticky_or_range362w364w & wire_w_lg_w_sticky_or_range359w361w & wire_w_lg_w_sticky_or_range356w358w & wire_w_lg_w_sticky_or_range353w355w & wire_w_lg_w_sticky_or_range350w352w & wire_w_lg_w_sticky_or_range347w349w & wire_w_lg_w_sticky_or_range344w346w & wire_w_lg_w_sticky_or_range341w343w & wire_w_lg_w_sticky_or_range338w340w & wire_w_lg_w_sticky_or_range335w337w & wire_w_lg_w_sticky_or_range332w334w & wire_w_lg_w_sticky_or_range329w331w & wire_w_lg_w_sticky_or_range326w328w & wire_w_lg_w_sticky_or_range323w325w & wire_w_lg_w_sticky_or_range320w322w & wire_w_lg_w_sticky_or_range317w319w & wire_w_lg_w_sticky_or_range314w316w & wire_w_lg_w_sticky_or_range311w313w & wire_w_lg_w_sticky_or_range308w310w & wire_w_lg_w_sticky_or_range305w307w & wire_w_lg_w_sticky_or_range302w304w & wire_w_lg_w_sticky_or_range299w301w & wire_w_lg_w_sticky_or_range296w298w & wire_w_lg_w_sticky_or_range293w295w & wire_w_lg_w_sticky_or_range290w292w & wire_w_lg_w_sticky_or_range286w289w & sticky_bus(0));
	unsigned_integer <= integer_rounded_reg;
	upper_limit_w <= ((wire_sign_input_reg3_w_lg_q458w(0) AND (exceed_upper_limit_reg3 OR equal_upper_limit_reg3)) OR wire_sign_input_reg3_w_lg_q456w(0));
	zero_input_w <= (wire_exp_or_reg4_w_lg_q220w(0) AND wire_man_or_reg4_w_lg_q222w(0));
	wire_w_below_lower_limit3_anding_range228w(0) <= below_lower_limit3_anding(0);
	wire_w_below_lower_limit3_anding_range232w(0) <= below_lower_limit3_anding(1);
	wire_w_below_lower_limit3_anding_range235w(0) <= below_lower_limit3_anding(2);
	wire_w_below_lower_limit3_anding_range238w(0) <= below_lower_limit3_anding(3);
	wire_w_below_lower_limit3_anding_range241w(0) <= below_lower_limit3_anding(4);
	wire_w_below_lower_limit3_anding_range244w(0) <= below_lower_limit3_anding(5);
	wire_w_below_lower_limit3_anding_range247w(0) <= below_lower_limit3_anding(6);
	wire_w_below_lower_limit3_anding_range250w(0) <= below_lower_limit3_anding(7);
	wire_w_below_lower_limit3_anding_range253w(0) <= below_lower_limit3_anding(8);
	wire_w_below_lower_limit3_anding_range256w(0) <= below_lower_limit3_anding(9);
	wire_w_below_lower_limit3_oring_range260w(0) <= below_lower_limit3_oring(0);
	wire_w_below_lower_limit3_oring_range263w(0) <= below_lower_limit3_oring(1);
	wire_w_below_lower_limit3_oring_range265w(0) <= below_lower_limit3_oring(2);
	wire_w_below_lower_limit3_oring_range267w(0) <= below_lower_limit3_oring(3);
	wire_w_exp_and_range8w(0) <= exp_and(0);
	wire_w_exp_and_range14w(0) <= exp_and(1);
	wire_w_exp_and_range19w(0) <= exp_and(2);
	wire_w_exp_and_range24w(0) <= exp_and(3);
	wire_w_exp_and_range29w(0) <= exp_and(4);
	wire_w_exp_and_range34w(0) <= exp_and(5);
	wire_w_exp_and_range39w(0) <= exp_and(6);
	wire_w_exp_and_range44w(0) <= exp_and(7);
	wire_w_exp_and_range49w(0) <= exp_and(8);
	wire_w_exp_and_range54w(0) <= exp_and(9);
	wire_w_exp_bus_range55w(0) <= exp_bus(10);
	wire_w_exp_bus_range10w(0) <= exp_bus(1);
	wire_w_exp_bus_range15w(0) <= exp_bus(2);
	wire_w_exp_bus_range20w(0) <= exp_bus(3);
	wire_w_exp_bus_range25w(0) <= exp_bus(4);
	wire_w_exp_bus_range30w(0) <= exp_bus(5);
	wire_w_exp_bus_range35w(0) <= exp_bus(6);
	wire_w_exp_bus_range40w(0) <= exp_bus(7);
	wire_w_exp_bus_range45w(0) <= exp_bus(8);
	wire_w_exp_bus_range50w(0) <= exp_bus(9);
	wire_w_exp_or_range6w(0) <= exp_or(0);
	wire_w_exp_or_range12w(0) <= exp_or(1);
	wire_w_exp_or_range17w(0) <= exp_or(2);
	wire_w_exp_or_range22w(0) <= exp_or(3);
	wire_w_exp_or_range27w(0) <= exp_or(4);
	wire_w_exp_or_range32w(0) <= exp_or(5);
	wire_w_exp_or_range37w(0) <= exp_or(6);
	wire_w_exp_or_range42w(0) <= exp_or(7);
	wire_w_exp_or_range47w(0) <= exp_or(8);
	wire_w_exp_or_range52w(0) <= exp_or(9);
	wire_w_inv_integer_range452w <= inv_integer(62 DOWNTO 31);
	wire_w_man_bus1_range136w(0) <= man_bus1(0);
	wire_w_man_bus1_range106w(0) <= man_bus1(10);
	wire_w_man_bus1_range103w(0) <= man_bus1(11);
	wire_w_man_bus1_range100w(0) <= man_bus1(12);
	wire_w_man_bus1_range97w(0) <= man_bus1(13);
	wire_w_man_bus1_range94w(0) <= man_bus1(14);
	wire_w_man_bus1_range91w(0) <= man_bus1(15);
	wire_w_man_bus1_range88w(0) <= man_bus1(16);
	wire_w_man_bus1_range85w(0) <= man_bus1(17);
	wire_w_man_bus1_range82w(0) <= man_bus1(18);
	wire_w_man_bus1_range79w(0) <= man_bus1(19);
	wire_w_man_bus1_range133w(0) <= man_bus1(1);
	wire_w_man_bus1_range76w(0) <= man_bus1(20);
	wire_w_man_bus1_range73w(0) <= man_bus1(21);
	wire_w_man_bus1_range70w(0) <= man_bus1(22);
	wire_w_man_bus1_range67w(0) <= man_bus1(23);
	wire_w_man_bus1_range64w(0) <= man_bus1(24);
	wire_w_man_bus1_range130w(0) <= man_bus1(2);
	wire_w_man_bus1_range127w(0) <= man_bus1(3);
	wire_w_man_bus1_range124w(0) <= man_bus1(4);
	wire_w_man_bus1_range121w(0) <= man_bus1(5);
	wire_w_man_bus1_range118w(0) <= man_bus1(6);
	wire_w_man_bus1_range115w(0) <= man_bus1(7);
	wire_w_man_bus1_range112w(0) <= man_bus1(8);
	wire_w_man_bus1_range109w(0) <= man_bus1(9);
	wire_w_man_bus2_range215w(0) <= man_bus2(0);
	wire_w_man_bus2_range185w(0) <= man_bus2(10);
	wire_w_man_bus2_range182w(0) <= man_bus2(11);
	wire_w_man_bus2_range179w(0) <= man_bus2(12);
	wire_w_man_bus2_range176w(0) <= man_bus2(13);
	wire_w_man_bus2_range173w(0) <= man_bus2(14);
	wire_w_man_bus2_range170w(0) <= man_bus2(15);
	wire_w_man_bus2_range167w(0) <= man_bus2(16);
	wire_w_man_bus2_range164w(0) <= man_bus2(17);
	wire_w_man_bus2_range161w(0) <= man_bus2(18);
	wire_w_man_bus2_range158w(0) <= man_bus2(19);
	wire_w_man_bus2_range212w(0) <= man_bus2(1);
	wire_w_man_bus2_range155w(0) <= man_bus2(20);
	wire_w_man_bus2_range152w(0) <= man_bus2(21);
	wire_w_man_bus2_range149w(0) <= man_bus2(22);
	wire_w_man_bus2_range146w(0) <= man_bus2(23);
	wire_w_man_bus2_range143w(0) <= man_bus2(24);
	wire_w_man_bus2_range209w(0) <= man_bus2(2);
	wire_w_man_bus2_range206w(0) <= man_bus2(3);
	wire_w_man_bus2_range203w(0) <= man_bus2(4);
	wire_w_man_bus2_range200w(0) <= man_bus2(5);
	wire_w_man_bus2_range197w(0) <= man_bus2(6);
	wire_w_man_bus2_range194w(0) <= man_bus2(7);
	wire_w_man_bus2_range191w(0) <= man_bus2(8);
	wire_w_man_bus2_range188w(0) <= man_bus2(9);
	wire_w_man_or1_range108w(0) <= man_or1(10);
	wire_w_man_or1_range105w(0) <= man_or1(11);
	wire_w_man_or1_range102w(0) <= man_or1(12);
	wire_w_man_or1_range99w(0) <= man_or1(13);
	wire_w_man_or1_range96w(0) <= man_or1(14);
	wire_w_man_or1_range93w(0) <= man_or1(15);
	wire_w_man_or1_range90w(0) <= man_or1(16);
	wire_w_man_or1_range87w(0) <= man_or1(17);
	wire_w_man_or1_range84w(0) <= man_or1(18);
	wire_w_man_or1_range81w(0) <= man_or1(19);
	wire_w_man_or1_range135w(0) <= man_or1(1);
	wire_w_man_or1_range78w(0) <= man_or1(20);
	wire_w_man_or1_range75w(0) <= man_or1(21);
	wire_w_man_or1_range72w(0) <= man_or1(22);
	wire_w_man_or1_range69w(0) <= man_or1(23);
	wire_w_man_or1_range66w(0) <= man_or1(24);
	wire_w_man_or1_range62w(0) <= man_or1(25);
	wire_w_man_or1_range132w(0) <= man_or1(2);
	wire_w_man_or1_range129w(0) <= man_or1(3);
	wire_w_man_or1_range126w(0) <= man_or1(4);
	wire_w_man_or1_range123w(0) <= man_or1(5);
	wire_w_man_or1_range120w(0) <= man_or1(6);
	wire_w_man_or1_range117w(0) <= man_or1(7);
	wire_w_man_or1_range114w(0) <= man_or1(8);
	wire_w_man_or1_range111w(0) <= man_or1(9);
	wire_w_man_or2_range187w(0) <= man_or2(10);
	wire_w_man_or2_range184w(0) <= man_or2(11);
	wire_w_man_or2_range181w(0) <= man_or2(12);
	wire_w_man_or2_range178w(0) <= man_or2(13);
	wire_w_man_or2_range175w(0) <= man_or2(14);
	wire_w_man_or2_range172w(0) <= man_or2(15);
	wire_w_man_or2_range169w(0) <= man_or2(16);
	wire_w_man_or2_range166w(0) <= man_or2(17);
	wire_w_man_or2_range163w(0) <= man_or2(18);
	wire_w_man_or2_range160w(0) <= man_or2(19);
	wire_w_man_or2_range214w(0) <= man_or2(1);
	wire_w_man_or2_range157w(0) <= man_or2(20);
	wire_w_man_or2_range154w(0) <= man_or2(21);
	wire_w_man_or2_range151w(0) <= man_or2(22);
	wire_w_man_or2_range148w(0) <= man_or2(23);
	wire_w_man_or2_range145w(0) <= man_or2(24);
	wire_w_man_or2_range141w(0) <= man_or2(25);
	wire_w_man_or2_range211w(0) <= man_or2(2);
	wire_w_man_or2_range208w(0) <= man_or2(3);
	wire_w_man_or2_range205w(0) <= man_or2(4);
	wire_w_man_or2_range202w(0) <= man_or2(5);
	wire_w_man_or2_range199w(0) <= man_or2(6);
	wire_w_man_or2_range196w(0) <= man_or2(7);
	wire_w_man_or2_range193w(0) <= man_or2(8);
	wire_w_man_or2_range190w(0) <= man_or2(9);
	wire_w_sticky_bus_range315w(0) <= sticky_bus(10);
	wire_w_sticky_bus_range318w(0) <= sticky_bus(11);
	wire_w_sticky_bus_range321w(0) <= sticky_bus(12);
	wire_w_sticky_bus_range324w(0) <= sticky_bus(13);
	wire_w_sticky_bus_range327w(0) <= sticky_bus(14);
	wire_w_sticky_bus_range330w(0) <= sticky_bus(15);
	wire_w_sticky_bus_range333w(0) <= sticky_bus(16);
	wire_w_sticky_bus_range336w(0) <= sticky_bus(17);
	wire_w_sticky_bus_range339w(0) <= sticky_bus(18);
	wire_w_sticky_bus_range342w(0) <= sticky_bus(19);
	wire_w_sticky_bus_range288w(0) <= sticky_bus(1);
	wire_w_sticky_bus_range345w(0) <= sticky_bus(20);
	wire_w_sticky_bus_range348w(0) <= sticky_bus(21);
	wire_w_sticky_bus_range351w(0) <= sticky_bus(22);
	wire_w_sticky_bus_range354w(0) <= sticky_bus(23);
	wire_w_sticky_bus_range357w(0) <= sticky_bus(24);
	wire_w_sticky_bus_range360w(0) <= sticky_bus(25);
	wire_w_sticky_bus_range363w(0) <= sticky_bus(26);
	wire_w_sticky_bus_range366w(0) <= sticky_bus(27);
	wire_w_sticky_bus_range369w(0) <= sticky_bus(28);
	wire_w_sticky_bus_range372w(0) <= sticky_bus(29);
	wire_w_sticky_bus_range291w(0) <= sticky_bus(2);
	wire_w_sticky_bus_range375w(0) <= sticky_bus(30);
	wire_w_sticky_bus_range378w(0) <= sticky_bus(31);
	wire_w_sticky_bus_range381w(0) <= sticky_bus(32);
	wire_w_sticky_bus_range384w(0) <= sticky_bus(33);
	wire_w_sticky_bus_range387w(0) <= sticky_bus(34);
	wire_w_sticky_bus_range390w(0) <= sticky_bus(35);
	wire_w_sticky_bus_range393w(0) <= sticky_bus(36);
	wire_w_sticky_bus_range396w(0) <= sticky_bus(37);
	wire_w_sticky_bus_range399w(0) <= sticky_bus(38);
	wire_w_sticky_bus_range402w(0) <= sticky_bus(39);
	wire_w_sticky_bus_range294w(0) <= sticky_bus(3);
	wire_w_sticky_bus_range405w(0) <= sticky_bus(40);
	wire_w_sticky_bus_range408w(0) <= sticky_bus(41);
	wire_w_sticky_bus_range411w(0) <= sticky_bus(42);
	wire_w_sticky_bus_range414w(0) <= sticky_bus(43);
	wire_w_sticky_bus_range417w(0) <= sticky_bus(44);
	wire_w_sticky_bus_range420w(0) <= sticky_bus(45);
	wire_w_sticky_bus_range423w(0) <= sticky_bus(46);
	wire_w_sticky_bus_range426w(0) <= sticky_bus(47);
	wire_w_sticky_bus_range429w(0) <= sticky_bus(48);
	wire_w_sticky_bus_range432w(0) <= sticky_bus(49);
	wire_w_sticky_bus_range297w(0) <= sticky_bus(4);
	wire_w_sticky_bus_range435w(0) <= sticky_bus(50);
	wire_w_sticky_bus_range300w(0) <= sticky_bus(5);
	wire_w_sticky_bus_range303w(0) <= sticky_bus(6);
	wire_w_sticky_bus_range306w(0) <= sticky_bus(7);
	wire_w_sticky_bus_range309w(0) <= sticky_bus(8);
	wire_w_sticky_bus_range312w(0) <= sticky_bus(9);
	wire_w_sticky_or_range286w(0) <= sticky_or(0);
	wire_w_sticky_or_range317w(0) <= sticky_or(10);
	wire_w_sticky_or_range320w(0) <= sticky_or(11);
	wire_w_sticky_or_range323w(0) <= sticky_or(12);
	wire_w_sticky_or_range326w(0) <= sticky_or(13);
	wire_w_sticky_or_range329w(0) <= sticky_or(14);
	wire_w_sticky_or_range332w(0) <= sticky_or(15);
	wire_w_sticky_or_range335w(0) <= sticky_or(16);
	wire_w_sticky_or_range338w(0) <= sticky_or(17);
	wire_w_sticky_or_range341w(0) <= sticky_or(18);
	wire_w_sticky_or_range344w(0) <= sticky_or(19);
	wire_w_sticky_or_range290w(0) <= sticky_or(1);
	wire_w_sticky_or_range347w(0) <= sticky_or(20);
	wire_w_sticky_or_range350w(0) <= sticky_or(21);
	wire_w_sticky_or_range353w(0) <= sticky_or(22);
	wire_w_sticky_or_range356w(0) <= sticky_or(23);
	wire_w_sticky_or_range359w(0) <= sticky_or(24);
	wire_w_sticky_or_range362w(0) <= sticky_or(25);
	wire_w_sticky_or_range365w(0) <= sticky_or(26);
	wire_w_sticky_or_range368w(0) <= sticky_or(27);
	wire_w_sticky_or_range371w(0) <= sticky_or(28);
	wire_w_sticky_or_range374w(0) <= sticky_or(29);
	wire_w_sticky_or_range293w(0) <= sticky_or(2);
	wire_w_sticky_or_range377w(0) <= sticky_or(30);
	wire_w_sticky_or_range380w(0) <= sticky_or(31);
	wire_w_sticky_or_range383w(0) <= sticky_or(32);
	wire_w_sticky_or_range386w(0) <= sticky_or(33);
	wire_w_sticky_or_range389w(0) <= sticky_or(34);
	wire_w_sticky_or_range392w(0) <= sticky_or(35);
	wire_w_sticky_or_range395w(0) <= sticky_or(36);
	wire_w_sticky_or_range398w(0) <= sticky_or(37);
	wire_w_sticky_or_range401w(0) <= sticky_or(38);
	wire_w_sticky_or_range404w(0) <= sticky_or(39);
	wire_w_sticky_or_range296w(0) <= sticky_or(3);
	wire_w_sticky_or_range407w(0) <= sticky_or(40);
	wire_w_sticky_or_range410w(0) <= sticky_or(41);
	wire_w_sticky_or_range413w(0) <= sticky_or(42);
	wire_w_sticky_or_range416w(0) <= sticky_or(43);
	wire_w_sticky_or_range419w(0) <= sticky_or(44);
	wire_w_sticky_or_range422w(0) <= sticky_or(45);
	wire_w_sticky_or_range425w(0) <= sticky_or(46);
	wire_w_sticky_or_range428w(0) <= sticky_or(47);
	wire_w_sticky_or_range431w(0) <= sticky_or(48);
	wire_w_sticky_or_range434w(0) <= sticky_or(49);
	wire_w_sticky_or_range299w(0) <= sticky_or(4);
	wire_w_sticky_or_range302w(0) <= sticky_or(5);
	wire_w_sticky_or_range305w(0) <= sticky_or(6);
	wire_w_sticky_or_range308w(0) <= sticky_or(7);
	wire_w_sticky_or_range311w(0) <= sticky_or(8);
	wire_w_sticky_or_range314w(0) <= sticky_or(9);
	wire_altbarrel_shift2_distance <= wire_w_lg_w_lg_barrel_direction_negative279w280w;
	loop49 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_barrel_direction_negative279w280w(i) <= wire_w_lg_barrel_direction_negative279w(i) OR wire_w_lg_w_lg_barrel_direction_negative277w278w(i);
	END GENERATE loop49;
	altbarrel_shift2 :  tofixed_altbarrel_shift_v5h
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => barrel_mantissa_input,
		direction => barrel_direction_negative,
		distance => wire_altbarrel_shift2_distance,
		result => wire_altbarrel_shift2_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN added_power2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN added_power2_reg <= wire_add_sub1_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_direction_negative_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_direction_negative_reg <= wire_power2_value_w_result_range257w(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg1 <= below_lower_limit3_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg2 <= below_lower_limit3_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg3 <= below_lower_limit3_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit3_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit3_reg4 <= below_lower_limit3_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg1 <= wire_below_lower_limit2_aeb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg2 <= border_lower_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg3 <= border_lower_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN border_lower_limit_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN border_lower_limit_reg4 <= border_lower_limit_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_border_lower_limit_reg4_w_lg_q489w(0) <= NOT border_lower_limit_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_reg <= dataa;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg1 <= equal_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg2 <= equal_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg3 <= equal_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_equal_upper_limit_reg3_w_lg_q454w(0) <= equal_upper_limit_reg3 AND wire_int_or_reg3_w_lg_q453w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg1 <= exceed_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg2 <= exceed_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg3 <= exceed_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_exceed_upper_limit_reg3_w_lg_q455w(0) <= exceed_upper_limit_reg3 OR wire_equal_upper_limit_reg3_w_lg_q454w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg4 <= upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg1 <= exp_and_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg2 <= exp_and_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg3 <= exp_and_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg4 <= exp_and_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg1 <= exp_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg2 <= exp_or_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg3 <= exp_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg4 <= exp_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_or_reg4_w_lg_q220w(0) <= NOT exp_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or1_reg1 <= int_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or2_reg1 <= int_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg2 <= (int_or1_reg1 OR int_or2_reg1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg3 <= int_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_int_or_reg3_w_lg_q453w(0) <= int_or_reg3 OR add_1_w;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_result_reg <= integer_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_rounded_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_rounded_reg <= integer_rounded;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or1_reg1 <= man_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or2_reg1 <= man_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg2 <= man_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg3 <= man_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg4 <= man_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_man_or_reg4_w_lg_q222w(0) <= NOT man_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_input_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_input_reg <= mantissa_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_exceeder_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_exceeder_reg <= more_than_max_shift_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_reg <= wire_max_shift_compare_agb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN power2_value_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN power2_value_reg <= power2_value_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg1 <= sign_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg2 <= sign_input_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg3 <= sign_input_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_input_reg3_w_lg_q456w(0) <= sign_input_reg3 AND wire_exceed_upper_limit_reg3_w_lg_q455w(0);
	wire_sign_input_reg3_w_lg_q458w(0) <= NOT sign_input_reg3;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg4 <= sign_input_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_add_1_adder_datab <= "000000000000000000000000000000000000000000000000000000000000001";
	add_1_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 63,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_1_adder_cout,
		dataa => integer_pre_round,
		datab => wire_add_1_adder_datab,
		result => wire_add_1_adder_result
	  );
	wire_add_sub1_datab <= "0000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 7,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => power2_value_reg,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	loop50 : FOR i IN 0 TO 31 GENERATE 
		wire_add_sub3_w_lg_w_lg_cout465w466w(i) <= wire_add_sub3_w_lg_cout465w(0) AND wire_w_inv_integer_range452w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 31 GENERATE 
		wire_add_sub3_w_lg_cout464w(i) <= wire_add_sub3_cout AND wire_add_sub4_result(i);
	END GENERATE loop51;
	wire_add_sub3_w_lg_cout465w(0) <= NOT wire_add_sub3_cout;
	wire_add_sub3_datab <= "0000000000000000000000000000001";
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 31,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub3_cout,
		dataa => inv_integer(30 DOWNTO 0),
		datab => wire_add_sub3_datab,
		result => wire_add_sub3_result
	  );
	wire_add_sub4_datab <= "00000000000000000000000000000001";
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 32,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => inv_integer(62 DOWNTO 31),
		datab => wire_add_sub4_datab,
		result => wire_add_sub4_result
	  );
	wire_barrel_direction_invert_dataa <= (OTHERS => '0');
	barrel_direction_invert :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 7,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => wire_barrel_direction_invert_dataa,
		datab => power2_value_reg,
		result => wire_barrel_direction_invert_result
	  );
	wire_power2_value_w_lg_w_result_range257w269w(0) <= wire_power2_value_w_result_range257w(0) AND wire_w_below_lower_limit3_oring_range267w(0);
	wire_power2_value_w_lg_w_lg_w_result_range257w269w270w(0) <= wire_power2_value_w_lg_w_result_range257w269w(0) OR power2_value_overflow_w;
	wire_power2_value_w_result_range257w(0) <= wire_power2_value_result(10);
	wire_power2_value_w_result_range230w(0) <= wire_power2_value_result(1);
	wire_power2_value_w_result_range233w(0) <= wire_power2_value_result(2);
	wire_power2_value_w_result_range236w(0) <= wire_power2_value_result(3);
	wire_power2_value_w_result_range239w(0) <= wire_power2_value_result(4);
	wire_power2_value_w_result_range242w(0) <= wire_power2_value_result(5);
	wire_power2_value_w_result_range245w(0) <= wire_power2_value_result(6);
	wire_power2_value_w_result_range248w(0) <= wire_power2_value_result(7);
	wire_power2_value_w_result_range251w(0) <= wire_power2_value_result(8);
	wire_power2_value_w_result_range254w(0) <= wire_power2_value_result(9);
	power2_value :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_input,
		datab => shift_value_w,
		overflow => wire_power2_value_overflow,
		result => wire_power2_value_result
	  );
	below_lower_limit1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		aeb => wire_below_lower_limit1_aeb,
		dataa => exponent_input,
		datab => bias_value_less_1_w
	  );
	below_lower_limit2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		aeb => wire_below_lower_limit2_aeb,
		dataa => exponent_input,
		datab => shift_value_w
	  );
	exceed_upper_limit :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		aeb => wire_exceed_upper_limit_aeb,
		agb => wire_exceed_upper_limit_agb,
		dataa => padded_exponent_input,
		datab => const_bias_value_add_width_res_w
	  );
	max_shift_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 7
	  )
	  PORT MAP ( 
		agb => wire_max_shift_compare_agb,
		dataa => added_power2_reg,
		datab => max_shift_w
	  );

 END RTL; --tofixed_altfp_convert_2gn
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY tofixed IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END tofixed;


ARCHITECTURE RTL OF tofixed IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (63 DOWNTO 0);



	COMPONENT tofixed_altfp_convert_2gn
	PORT (
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(63 DOWNTO 0);

	tofixed_altfp_convert_2gn_component : tofixed_altfp_convert_2gn
	PORT MAP (
		aclr => aclr,
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "FLOAT2FIXED"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "64"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "11"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "12"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "52"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "64"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 64 0 INPUT NODEFVAL "dataa[63..0]"
-- Retrieval info: CONNECT: @dataa 0 0 64 0 dataa 0 0 64 0
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL tofixed.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL tofixed.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL tofixed.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL tofixed_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL tofixed.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL tofixed.cmp TRUE TRUE
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX NUMERIC "1"
-- Retrieval info: LIB_FILE: lpm
