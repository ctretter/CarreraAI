﻿-------------------------------------------------------------------------------
-- Title      : <Short title for this unit>
-- Project    : <Name of the design project>
-------------------------------------------------------------------------------
-- RevCtrl    : $Id: Template-e.vhd 63 2011-11-05 14:02:00Z mroland $
-- Author     : <Author(s) of this file>
-------------------------------------------------------------------------------
-- Description: <Detailed description of this unit's purpose>
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.global.all;

entity Template is
  
  generic (
    -- Your generics here
  );
  
  port (
    iClk         : in  std_ulogic;
    inResetAsync : in  std_ulogic;

    -- Your ports here
  );

end Template;
