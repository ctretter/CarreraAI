-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: FloatConv.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.0.0 Build 211 04/27/2016 SJ Standard Edition
-- ************************************************************


--Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="FIXED2FLOAT" ROUNDING="TO_NEAREST" WIDTH_DATA=64 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=11 WIDTH_INT=12 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=52 WIDTH_RESULT=64 aclr clock dataa result
--VERSION_BEGIN 16.0 cbx_altbarrel_shift 2016:04:27:18:05:34:SJ cbx_altera_syncram_nd_impl 2016:04:27:18:05:34:SJ cbx_altfp_convert 2016:04:27:18:05:34:SJ cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_altsyncram 2016:04:27:18:05:34:SJ cbx_cycloneii 2016:04:27:18:05:34:SJ cbx_lpm_abs 2016:04:27:18:05:34:SJ cbx_lpm_add_sub 2016:04:27:18:05:34:SJ cbx_lpm_compare 2016:04:27:18:05:34:SJ cbx_lpm_decode 2016:04:27:18:05:34:SJ cbx_lpm_divide 2016:04:27:18:05:34:SJ cbx_lpm_mux 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ cbx_nadder 2016:04:27:18:05:34:SJ cbx_stratix 2016:04:27:18:05:34:SJ cbx_stratixii 2016:04:27:18:05:34:SJ cbx_stratixiii 2016:04:27:18:05:34:SJ cbx_stratixv 2016:04:27:18:05:34:SJ cbx_util_mgl 2016:04:27:18:05:34:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=64 WIDTHDIST=6 aclr clk_en clock data distance result
--VERSION_BEGIN 16.0 cbx_altbarrel_shift 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END

--synthesis_resources = reg 133 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altbarrel_shift_lof IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END FloatConv_altbarrel_shift_lof;

 ARCHITECTURE RTL OF FloatConv_altbarrel_shift_lof IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec5r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w106w107w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w102w103w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w127w128w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w123w124w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w149w150w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w145w146w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w171w172w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w167w168w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w190w191w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w186w187w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w211w212w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w207w208w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w98w99w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w119w120w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w141w142w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w163w164w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w182w183w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w203w204w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range94w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range94w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range115w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range115w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range137w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range137w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range160w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range160w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range179w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range179w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range200w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range200w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_dir_w_range91w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_dir_w_range113w126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_dir_w_range134w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_dir_w_range158w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_dir_w_range177w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_dir_w_range197w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range94w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range115w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range137w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range160w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range179w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_sel_w_range200w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range94w106w107w108w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range115w127w128w129w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range137w149w150w151w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range160w171w172w173w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range179w190w191w192w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range200w211w212w213w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w109w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w130w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w152w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w174w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w193w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w214w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (447 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (383 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w101w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w104w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w122w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w125w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w144w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w147w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w166w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w169w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w185w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w188w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w206w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w209w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_dir_w_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_dir_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_dir_w_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_dir_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_dir_w_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_dir_w_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sbit_w_range112w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sbit_w_range132w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sbit_w_range154w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sbit_w_range176w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sbit_w_range195w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sbit_w_range89w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sel_w_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sel_w_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sel_w_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sel_w_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sel_w_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_sel_w_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_smux_w_range153w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_w_smux_w_range215w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w106w107w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range94w106w(0) AND wire_altbarrel_shift3_w104w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w102w103w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range94w102w(0) AND wire_altbarrel_shift3_w101w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w127w128w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range115w127w(0) AND wire_altbarrel_shift3_w125w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w123w124w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range115w123w(0) AND wire_altbarrel_shift3_w122w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w149w150w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range137w149w(0) AND wire_altbarrel_shift3_w147w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w145w146w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range137w145w(0) AND wire_altbarrel_shift3_w144w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w171w172w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range160w171w(0) AND wire_altbarrel_shift3_w169w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w167w168w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range160w167w(0) AND wire_altbarrel_shift3_w166w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w190w191w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range179w190w(0) AND wire_altbarrel_shift3_w188w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w186w187w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range179w186w(0) AND wire_altbarrel_shift3_w185w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w211w212w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range200w211w(0) AND wire_altbarrel_shift3_w209w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w207w208w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range200w207w(0) AND wire_altbarrel_shift3_w206w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w98w99w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range94w98w(0) AND wire_altbarrel_shift3_w_sbit_w_range89w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w119w120w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range115w119w(0) AND wire_altbarrel_shift3_w_sbit_w_range112w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w141w142w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range137w141w(0) AND wire_altbarrel_shift3_w_sbit_w_range132w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w163w164w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range160w163w(0) AND wire_altbarrel_shift3_w_sbit_w_range154w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w182w183w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range179w182w(0) AND wire_altbarrel_shift3_w_sbit_w_range176w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w203w204w(i) <= wire_altbarrel_shift3_w_lg_w_sel_w_range200w203w(0) AND wire_altbarrel_shift3_w_sbit_w_range195w(i);
	END GENERATE loop17;
	wire_altbarrel_shift3_w_lg_w_sel_w_range94w106w(0) <= wire_altbarrel_shift3_w_sel_w_range94w(0) AND wire_altbarrel_shift3_w_lg_w_dir_w_range91w105w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range94w102w(0) <= wire_altbarrel_shift3_w_sel_w_range94w(0) AND wire_altbarrel_shift3_w_dir_w_range91w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range115w127w(0) <= wire_altbarrel_shift3_w_sel_w_range115w(0) AND wire_altbarrel_shift3_w_lg_w_dir_w_range113w126w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range115w123w(0) <= wire_altbarrel_shift3_w_sel_w_range115w(0) AND wire_altbarrel_shift3_w_dir_w_range113w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range137w149w(0) <= wire_altbarrel_shift3_w_sel_w_range137w(0) AND wire_altbarrel_shift3_w_lg_w_dir_w_range134w148w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range137w145w(0) <= wire_altbarrel_shift3_w_sel_w_range137w(0) AND wire_altbarrel_shift3_w_dir_w_range134w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range160w171w(0) <= wire_altbarrel_shift3_w_sel_w_range160w(0) AND wire_altbarrel_shift3_w_lg_w_dir_w_range158w170w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range160w167w(0) <= wire_altbarrel_shift3_w_sel_w_range160w(0) AND wire_altbarrel_shift3_w_dir_w_range158w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range179w190w(0) <= wire_altbarrel_shift3_w_sel_w_range179w(0) AND wire_altbarrel_shift3_w_lg_w_dir_w_range177w189w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range179w186w(0) <= wire_altbarrel_shift3_w_sel_w_range179w(0) AND wire_altbarrel_shift3_w_dir_w_range177w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range200w211w(0) <= wire_altbarrel_shift3_w_sel_w_range200w(0) AND wire_altbarrel_shift3_w_lg_w_dir_w_range197w210w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range200w207w(0) <= wire_altbarrel_shift3_w_sel_w_range200w(0) AND wire_altbarrel_shift3_w_dir_w_range197w(0);
	wire_altbarrel_shift3_w_lg_w_dir_w_range91w105w(0) <= NOT wire_altbarrel_shift3_w_dir_w_range91w(0);
	wire_altbarrel_shift3_w_lg_w_dir_w_range113w126w(0) <= NOT wire_altbarrel_shift3_w_dir_w_range113w(0);
	wire_altbarrel_shift3_w_lg_w_dir_w_range134w148w(0) <= NOT wire_altbarrel_shift3_w_dir_w_range134w(0);
	wire_altbarrel_shift3_w_lg_w_dir_w_range158w170w(0) <= NOT wire_altbarrel_shift3_w_dir_w_range158w(0);
	wire_altbarrel_shift3_w_lg_w_dir_w_range177w189w(0) <= NOT wire_altbarrel_shift3_w_dir_w_range177w(0);
	wire_altbarrel_shift3_w_lg_w_dir_w_range197w210w(0) <= NOT wire_altbarrel_shift3_w_dir_w_range197w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range94w98w(0) <= NOT wire_altbarrel_shift3_w_sel_w_range94w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range115w119w(0) <= NOT wire_altbarrel_shift3_w_sel_w_range115w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range137w141w(0) <= NOT wire_altbarrel_shift3_w_sel_w_range137w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range160w163w(0) <= NOT wire_altbarrel_shift3_w_sel_w_range160w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range179w182w(0) <= NOT wire_altbarrel_shift3_w_sel_w_range179w(0);
	wire_altbarrel_shift3_w_lg_w_sel_w_range200w203w(0) <= NOT wire_altbarrel_shift3_w_sel_w_range200w(0);
	loop18 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range94w106w107w108w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w106w107w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w102w103w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range115w127w128w129w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w127w128w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w123w124w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range137w149w150w151w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w149w150w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w145w146w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range160w171w172w173w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w171w172w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w167w168w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range179w190w191w192w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w190w191w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w186w187w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range200w211w212w213w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w211w212w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w207w208w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w109w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range94w106w107w108w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range94w98w99w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w130w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range115w127w128w129w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range115w119w120w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w152w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range137w149w150w151w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range137w141w142w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w174w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range160w171w172w173w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range160w163w164w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w193w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range179w190w191w192w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range179w182w183w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 63 GENERATE 
		wire_altbarrel_shift3_w214w(i) <= wire_altbarrel_shift3_w_lg_w_lg_w_lg_w_sel_w_range200w211w212w213w(i) OR wire_altbarrel_shift3_w_lg_w_lg_w_sel_w_range200w203w204w(i);
	END GENERATE loop29;
	dir_w <= ( dir_pipe(1) & dir_w(4 DOWNTO 3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(447 DOWNTO 384);
	sbit_w <= ( sbit_piper2d & smux_w(319 DOWNTO 192) & sbit_piper1d & smux_w(127 DOWNTO 0) & data);
	sel_w <= ( sel_pipec5r1d & sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift3_w214w & wire_altbarrel_shift3_w193w & wire_altbarrel_shift3_w174w & wire_altbarrel_shift3_w152w & wire_altbarrel_shift3_w130w & wire_altbarrel_shift3_w109w);
	wire_altbarrel_shift3_w101w <= ( pad_w(0) & sbit_w(63 DOWNTO 1));
	wire_altbarrel_shift3_w104w <= ( sbit_w(62 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift3_w122w <= ( pad_w(1 DOWNTO 0) & sbit_w(127 DOWNTO 66));
	wire_altbarrel_shift3_w125w <= ( sbit_w(125 DOWNTO 64) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift3_w144w <= ( pad_w(3 DOWNTO 0) & sbit_w(191 DOWNTO 132));
	wire_altbarrel_shift3_w147w <= ( sbit_w(187 DOWNTO 128) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift3_w166w <= ( pad_w(7 DOWNTO 0) & sbit_w(255 DOWNTO 200));
	wire_altbarrel_shift3_w169w <= ( sbit_w(247 DOWNTO 192) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift3_w185w <= ( pad_w(15 DOWNTO 0) & sbit_w(319 DOWNTO 272));
	wire_altbarrel_shift3_w188w <= ( sbit_w(303 DOWNTO 256) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift3_w206w <= ( pad_w(31 DOWNTO 0) & sbit_w(383 DOWNTO 352));
	wire_altbarrel_shift3_w209w <= ( sbit_w(351 DOWNTO 320) & pad_w(31 DOWNTO 0));
	wire_altbarrel_shift3_w_dir_w_range91w(0) <= dir_w(0);
	wire_altbarrel_shift3_w_dir_w_range113w(0) <= dir_w(1);
	wire_altbarrel_shift3_w_dir_w_range134w(0) <= dir_w(2);
	wire_altbarrel_shift3_w_dir_w_range158w(0) <= dir_w(3);
	wire_altbarrel_shift3_w_dir_w_range177w(0) <= dir_w(4);
	wire_altbarrel_shift3_w_dir_w_range197w(0) <= dir_w(5);
	wire_altbarrel_shift3_w_sbit_w_range112w <= sbit_w(127 DOWNTO 64);
	wire_altbarrel_shift3_w_sbit_w_range132w <= sbit_w(191 DOWNTO 128);
	wire_altbarrel_shift3_w_sbit_w_range154w <= sbit_w(255 DOWNTO 192);
	wire_altbarrel_shift3_w_sbit_w_range176w <= sbit_w(319 DOWNTO 256);
	wire_altbarrel_shift3_w_sbit_w_range195w <= sbit_w(383 DOWNTO 320);
	wire_altbarrel_shift3_w_sbit_w_range89w <= sbit_w(63 DOWNTO 0);
	wire_altbarrel_shift3_w_sel_w_range94w(0) <= sel_w(0);
	wire_altbarrel_shift3_w_sel_w_range115w(0) <= sel_w(1);
	wire_altbarrel_shift3_w_sel_w_range137w(0) <= sel_w(2);
	wire_altbarrel_shift3_w_sel_w_range160w(0) <= sel_w(3);
	wire_altbarrel_shift3_w_sel_w_range179w(0) <= sel_w(4);
	wire_altbarrel_shift3_w_sel_w_range200w(0) <= sel_w(5);
	wire_altbarrel_shift3_w_smux_w_range153w <= smux_w(191 DOWNTO 128);
	wire_altbarrel_shift3_w_smux_w_range215w <= smux_w(383 DOWNTO 320);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(5) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift3_w_smux_w_range153w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift3_w_smux_w_range215w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec5r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec5r1d <= distance(5);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --FloatConv_altbarrel_shift_lof


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=64 WIDTHAD=6 data q
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FloatConv_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --FloatConv_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FloatConv_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero260w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero262w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero260w & wire_altpriority_encoder16_w_lg_w_lg_zero262w263w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  FloatConv_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	wire_altpriority_encoder16_w_lg_w_lg_zero260w261w(0) <= wire_altpriority_encoder16_w_lg_zero260w(0) AND wire_altpriority_encoder16_q(0);
	wire_altpriority_encoder16_w_lg_zero262w(0) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(0);
	wire_altpriority_encoder16_w_lg_zero260w(0) <= NOT wire_altpriority_encoder16_zero;
	wire_altpriority_encoder16_w_lg_w_lg_zero262w263w(0) <= wire_altpriority_encoder16_w_lg_zero262w(0) OR wire_altpriority_encoder16_w_lg_w_lg_zero260w261w(0);
	altpriority_encoder16 :  FloatConv_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FloatConv_altpriority_encoder_be8;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero250w251w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero252w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero252w253w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero250w & wire_altpriority_encoder14_w_lg_w_lg_zero252w253w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  FloatConv_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop30 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero250w251w(i) <= wire_altpriority_encoder14_w_lg_zero250w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_zero252w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop31;
	wire_altpriority_encoder14_w_lg_zero250w(0) <= NOT wire_altpriority_encoder14_zero;
	loop32 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero252w253w(i) <= wire_altpriority_encoder14_w_lg_zero252w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero250w251w(i);
	END GENERATE loop32;
	altpriority_encoder14 :  FloatConv_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FloatConv_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero240w241w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero242w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero242w243w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero240w & wire_altpriority_encoder12_w_lg_w_lg_zero242w243w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  FloatConv_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	loop33 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero240w241w(i) <= wire_altpriority_encoder12_w_lg_zero240w(0) AND wire_altpriority_encoder12_q(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_zero242w(i) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(i);
	END GENERATE loop34;
	wire_altpriority_encoder12_w_lg_zero240w(0) <= NOT wire_altpriority_encoder12_zero;
	loop35 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero242w243w(i) <= wire_altpriority_encoder12_w_lg_zero242w(i) OR wire_altpriority_encoder12_w_lg_w_lg_zero240w241w(i);
	END GENERATE loop35;
	altpriority_encoder12 :  FloatConv_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_rf8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END FloatConv_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --FloatConv_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END FloatConv_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero294w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero296w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FloatConv_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero294w & wire_altpriority_encoder22_w_lg_w_lg_zero296w297w);
	altpriority_encoder21 :  FloatConv_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder21_q
	  );
	wire_altpriority_encoder22_w_lg_w_lg_zero294w295w(0) <= wire_altpriority_encoder22_w_lg_zero294w(0) AND wire_altpriority_encoder22_q(0);
	wire_altpriority_encoder22_w_lg_zero296w(0) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(0);
	wire_altpriority_encoder22_w_lg_zero294w(0) <= NOT wire_altpriority_encoder22_zero;
	wire_altpriority_encoder22_w_lg_w_lg_zero296w297w(0) <= wire_altpriority_encoder22_w_lg_zero296w(0) OR wire_altpriority_encoder22_w_lg_w_lg_zero294w295w(0);
	altpriority_encoder22 :  FloatConv_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_6v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END FloatConv_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero285w286w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero287w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero287w288w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FloatConv_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero285w & wire_altpriority_encoder20_w_lg_w_lg_zero287w288w);
	altpriority_encoder19 :  FloatConv_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop36 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero285w286w(i) <= wire_altpriority_encoder20_w_lg_zero285w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_zero287w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop37;
	wire_altpriority_encoder20_w_lg_zero285w(0) <= NOT wire_altpriority_encoder20_zero;
	loop38 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero287w288w(i) <= wire_altpriority_encoder20_w_lg_zero287w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero285w286w(i);
	END GENERATE loop38;
	altpriority_encoder20 :  FloatConv_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_bv7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END FloatConv_altpriority_encoder_r08;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero276w277w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero278w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero278w279w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FloatConv_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero276w & wire_altpriority_encoder18_w_lg_w_lg_zero278w279w);
	altpriority_encoder17 :  FloatConv_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	loop39 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero276w277w(i) <= wire_altpriority_encoder18_w_lg_zero276w(0) AND wire_altpriority_encoder18_q(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_zero278w(i) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(i);
	END GENERATE loop40;
	wire_altpriority_encoder18_w_lg_zero276w(0) <= NOT wire_altpriority_encoder18_zero;
	loop41 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero278w279w(i) <= wire_altpriority_encoder18_w_lg_zero278w(i) OR wire_altpriority_encoder18_w_lg_w_lg_zero276w277w(i);
	END GENERATE loop41;
	altpriority_encoder18 :  FloatConv_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_r08

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END FloatConv_altpriority_encoder_q08;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero231w232w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero233w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero233w234w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  FloatConv_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  FloatConv_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero231w & wire_altpriority_encoder10_w_lg_w_lg_zero233w234w);
	loop42 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero231w232w(i) <= wire_altpriority_encoder10_w_lg_zero231w(0) AND wire_altpriority_encoder10_q(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_zero233w(i) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(i);
	END GENERATE loop43;
	wire_altpriority_encoder10_w_lg_zero231w(0) <= NOT wire_altpriority_encoder10_zero;
	loop44 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero233w234w(i) <= wire_altpriority_encoder10_w_lg_zero233w(i) OR wire_altpriority_encoder10_w_lg_w_lg_zero231w232w(i);
	END GENERATE loop44;
	altpriority_encoder10 :  FloatConv_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  FloatConv_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --FloatConv_altpriority_encoder_q08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 16.0 cbx_altpriority_encoder 2016:04:27:18:05:34:SJ cbx_mgl 2016:04:27:18:06:48:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_qf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FloatConv_altpriority_encoder_qf8;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_qf8 IS

	 SIGNAL  wire_altpriority_encoder23_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder24_w_lg_w_lg_zero306w307w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_zero308w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_zero306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_w_lg_zero308w309w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder24_w_lg_zero306w & wire_altpriority_encoder24_w_lg_w_lg_zero308w309w);
	zero <= (wire_altpriority_encoder23_zero AND wire_altpriority_encoder24_zero);
	altpriority_encoder23 :  FloatConv_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder23_q,
		zero => wire_altpriority_encoder23_zero
	  );
	loop45 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder24_w_lg_w_lg_zero306w307w(i) <= wire_altpriority_encoder24_w_lg_zero306w(0) AND wire_altpriority_encoder24_q(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder24_w_lg_zero308w(i) <= wire_altpriority_encoder24_zero AND wire_altpriority_encoder23_q(i);
	END GENERATE loop46;
	wire_altpriority_encoder24_w_lg_zero306w(0) <= NOT wire_altpriority_encoder24_zero;
	loop47 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder24_w_lg_w_lg_zero308w309w(i) <= wire_altpriority_encoder24_w_lg_zero308w(i) OR wire_altpriority_encoder24_w_lg_w_lg_zero306w307w(i);
	END GENERATE loop47;
	altpriority_encoder24 :  FloatConv_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder24_q,
		zero => wire_altpriority_encoder24_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_qf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altpriority_encoder_0c6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END FloatConv_altpriority_encoder_0c6;

 ARCHITECTURE RTL OF FloatConv_altpriority_encoder_0c6 IS

	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero222w223w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero224w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero224w225w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_zero	:	STD_LOGIC;
	 COMPONENT  FloatConv_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FloatConv_altpriority_encoder_qf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder8_w_lg_zero222w & wire_altpriority_encoder8_w_lg_w_lg_zero224w225w);
	altpriority_encoder7 :  FloatConv_altpriority_encoder_q08
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder7_q
	  );
	loop48 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero222w223w(i) <= wire_altpriority_encoder8_w_lg_zero222w(0) AND wire_altpriority_encoder8_q(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder8_w_lg_zero224w(i) <= wire_altpriority_encoder8_zero AND wire_altpriority_encoder7_q(i);
	END GENERATE loop49;
	wire_altpriority_encoder8_w_lg_zero222w(0) <= NOT wire_altpriority_encoder8_zero;
	loop50 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero224w225w(i) <= wire_altpriority_encoder8_w_lg_zero224w(i) OR wire_altpriority_encoder8_w_lg_w_lg_zero222w223w(i);
	END GENERATE loop50;
	altpriority_encoder8 :  FloatConv_altpriority_encoder_qf8
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder8_q,
		zero => wire_altpriority_encoder8_zero
	  );

 END RTL; --FloatConv_altpriority_encoder_0c6

 LIBRARY lpm_ver;
 USE lpm_ver.all;

--synthesis_resources = lpm_add_sub 5 lpm_compare 1 reg 476 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FloatConv_altfp_convert_2gn IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END FloatConv_altfp_convert_2gn;

 ARCHITECTURE RTL OF FloatConv_altfp_convert_2gn IS

	 SIGNAL  wire_altbarrel_shift3_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift3_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL	 add_1_adder1_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_w_lg_q69w70w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q67w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_1_adder1_reg	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_reg	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_reg_w_lg_w_lg_q76w77w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q75w	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exponent_bus_pre_reg	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg2	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg3	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg	:	STD_LOGIC_VECTOR(62 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg2	:	STD_LOGIC_VECTOR(62 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissa_pre_round_reg	:	STD_LOGIC_VECTOR(52 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mantissa_pre_round_reg_w_q_range68w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL	 priority_encoder_reg	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_reg	:	STD_LOGIC_VECTOR(63 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_add_sub4_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub4_datab	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_add_sub5_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub5_datab	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_sub6_datab	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_exponent_value_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_below_bias_value_w_lg_w_lg_alb21w22w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_below_bias_value_w_lg_alb20w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_below_bias_value_w_lg_alb21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_below_bias_value_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_w61w62w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_w61w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mantissa_overflow80w81w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_max_neg_value_selector17w18w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_int_a5w6w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow79w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector16w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a4w	:	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range34w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range38w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range41w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range44w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range47w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range50w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range53w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range56w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_1_adder1_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  add_1_adder2_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  add_1_adder_w :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_int_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exceptions_value :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exponent_bus :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exponent_bus_pre :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exponent_output_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exponent_rounded :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exponent_zero_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  int_a :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  int_a_2s :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  invert_int_a :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  leading_zeroes :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mag_int_a :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  mantissa_bus :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  mantissa_overflow :	STD_LOGIC;
	 SIGNAL  mantissa_post_round :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  mantissa_pre_round :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  mantissa_rounded :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  max_neg_value_selector :	STD_LOGIC;
	 SIGNAL  max_neg_value_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  minus_leading_zero :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  prio_mag_int_a :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  shifted_mag_int_a :	STD_LOGIC_VECTOR (62 DOWNTO 0);
	 SIGNAL  sign_bus :	STD_LOGIC;
	 SIGNAL  sign_int_a :	STD_LOGIC;
	 SIGNAL  sticky_bit_bus :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  sticky_bit_or_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  zero_padding_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  FloatConv_altbarrel_shift_lof
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(63 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FloatConv_altpriority_encoder_0c6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_guard_bit_w61w62w63w(0) <= wire_w_lg_w_lg_guard_bit_w61w62w(0) AND sticky_bit_w;
	wire_w_lg_w_lg_guard_bit_w61w62w(0) <= wire_w_lg_guard_bit_w61w(0) AND round_bit_w;
	loop51 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_mantissa_overflow80w81w(i) <= wire_w_lg_mantissa_overflow80w(0) AND exponent_bus_pre_reg(i);
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_max_neg_value_selector17w18w(i) <= wire_w_lg_max_neg_value_selector17w(0) AND exponent_zero_w(i);
	END GENERATE loop52;
	loop53 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_w_lg_sign_int_a5w6w(i) <= wire_w_lg_sign_int_a5w(0) AND int_a(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_mantissa_overflow79w(i) <= mantissa_overflow AND wire_add_sub6_result(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_max_neg_value_selector16w(i) <= max_neg_value_selector AND max_neg_value_w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 62 GENERATE 
		wire_w_lg_sign_int_a4w(i) <= sign_int_a AND int_a_2s(i);
	END GENERATE loop56;
	wire_w_lg_guard_bit_w61w(0) <= NOT guard_bit_w;
	wire_w_lg_mantissa_overflow80w(0) <= NOT mantissa_overflow;
	wire_w_lg_max_neg_value_selector17w(0) <= NOT max_neg_value_selector;
	wire_w_lg_sign_int_a5w(0) <= NOT sign_int_a;
	wire_w_lg_w_sticky_bit_or_w_range34w37w(0) <= wire_w_sticky_bit_or_w_range34w(0) OR wire_w_sticky_bit_bus_range36w(0);
	wire_w_lg_w_sticky_bit_or_w_range38w40w(0) <= wire_w_sticky_bit_or_w_range38w(0) OR wire_w_sticky_bit_bus_range39w(0);
	wire_w_lg_w_sticky_bit_or_w_range41w43w(0) <= wire_w_sticky_bit_or_w_range41w(0) OR wire_w_sticky_bit_bus_range42w(0);
	wire_w_lg_w_sticky_bit_or_w_range44w46w(0) <= wire_w_sticky_bit_or_w_range44w(0) OR wire_w_sticky_bit_bus_range45w(0);
	wire_w_lg_w_sticky_bit_or_w_range47w49w(0) <= wire_w_sticky_bit_or_w_range47w(0) OR wire_w_sticky_bit_bus_range48w(0);
	wire_w_lg_w_sticky_bit_or_w_range50w52w(0) <= wire_w_sticky_bit_or_w_range50w(0) OR wire_w_sticky_bit_bus_range51w(0);
	wire_w_lg_w_sticky_bit_or_w_range53w55w(0) <= wire_w_sticky_bit_or_w_range53w(0) OR wire_w_sticky_bit_bus_range54w(0);
	wire_w_lg_w_sticky_bit_or_w_range56w58w(0) <= wire_w_sticky_bit_or_w_range56w(0) OR wire_w_sticky_bit_bus_range57w(0);
	add_1_adder1_w <= add_1_adder1_reg;
	add_1_adder2_w <= (wire_add_1_adder1_cout_reg_w_lg_w_lg_q69w70w OR wire_add_1_adder1_cout_reg_w_lg_q67w);
	add_1_adder_w <= ( add_1_adder2_w & add_1_adder1_w);
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_w61w62w63w(0) OR (guard_bit_w AND round_bit_w));
	bias_value_w <= "01111001011";
	clk_en <= '1';
	const_bias_value_add_width_int_w <= "10000001001";
	exceptions_value <= (wire_w_lg_w_lg_max_neg_value_selector17w18w OR wire_w_lg_max_neg_value_selector16w);
	exponent_bus <= exponent_rounded;
	exponent_bus_pre <= (wire_below_bias_value_w_lg_w_lg_alb21w22w OR wire_below_bias_value_w_lg_alb20w);
	exponent_output_w <= wire_exponent_value_result;
	exponent_rounded <= (wire_w_lg_w_lg_mantissa_overflow80w81w OR wire_w_lg_mantissa_overflow79w);
	exponent_zero_w <= (OTHERS => '0');
	guard_bit_w <= shifted_mag_int_a(10);
	int_a <= dataa(62 DOWNTO 0);
	int_a_2s <= wire_add_sub1_result;
	invert_int_a <= (NOT int_a);
	leading_zeroes <= (NOT priority_encoder_reg);
	mag_int_a <= (wire_w_lg_w_lg_sign_int_a5w6w OR wire_w_lg_sign_int_a4w);
	mantissa_bus <= mantissa_rounded(51 DOWNTO 0);
	mantissa_overflow <= ((add_1_reg AND add_1_adder1_cout_reg) AND add_1_adder2_cout_reg);
	mantissa_post_round <= add_1_adder_w;
	mantissa_pre_round <= shifted_mag_int_a(62 DOWNTO 10);
	mantissa_rounded <= (wire_add_1_reg_w_lg_w_lg_q76w77w OR wire_add_1_reg_w_lg_q75w);
	max_neg_value_selector <= (wire_below_bias_value_alb AND sign_int_a_reg2);
	max_neg_value_w <= "10000001010";
	minus_leading_zero <= ( zero_padding_w & leading_zeroes);
	prio_mag_int_a <= ( mag_int_a_reg & "1");
	result <= result_reg;
	result_w <= ( sign_bus & exponent_bus & mantissa_bus);
	round_bit_w <= shifted_mag_int_a(9);
	shifted_mag_int_a <= wire_altbarrel_shift3_result(62 DOWNTO 0);
	sign_bus <= sign_int_a_reg5;
	sign_int_a <= dataa(63);
	sticky_bit_bus <= shifted_mag_int_a(8 DOWNTO 0);
	sticky_bit_or_w <= ( wire_w_lg_w_sticky_bit_or_w_range56w58w & wire_w_lg_w_sticky_bit_or_w_range53w55w & wire_w_lg_w_sticky_bit_or_w_range50w52w & wire_w_lg_w_sticky_bit_or_w_range47w49w & wire_w_lg_w_sticky_bit_or_w_range44w46w & wire_w_lg_w_sticky_bit_or_w_range41w43w & wire_w_lg_w_sticky_bit_or_w_range38w40w & wire_w_lg_w_sticky_bit_or_w_range34w37w & sticky_bit_bus(0));
	sticky_bit_w <= sticky_bit_or_w(8);
	zero_padding_w <= (OTHERS => '0');
	wire_w_sticky_bit_bus_range36w(0) <= sticky_bit_bus(1);
	wire_w_sticky_bit_bus_range39w(0) <= sticky_bit_bus(2);
	wire_w_sticky_bit_bus_range42w(0) <= sticky_bit_bus(3);
	wire_w_sticky_bit_bus_range45w(0) <= sticky_bit_bus(4);
	wire_w_sticky_bit_bus_range48w(0) <= sticky_bit_bus(5);
	wire_w_sticky_bit_bus_range51w(0) <= sticky_bit_bus(6);
	wire_w_sticky_bit_bus_range54w(0) <= sticky_bit_bus(7);
	wire_w_sticky_bit_bus_range57w(0) <= sticky_bit_bus(8);
	wire_w_sticky_bit_or_w_range34w(0) <= sticky_bit_or_w(0);
	wire_w_sticky_bit_or_w_range38w(0) <= sticky_bit_or_w(1);
	wire_w_sticky_bit_or_w_range41w(0) <= sticky_bit_or_w(2);
	wire_w_sticky_bit_or_w_range44w(0) <= sticky_bit_or_w(3);
	wire_w_sticky_bit_or_w_range47w(0) <= sticky_bit_or_w(4);
	wire_w_sticky_bit_or_w_range50w(0) <= sticky_bit_or_w(5);
	wire_w_sticky_bit_or_w_range53w(0) <= sticky_bit_or_w(6);
	wire_w_sticky_bit_or_w_range56w(0) <= sticky_bit_or_w(7);
	wire_altbarrel_shift3_data <= ( "0" & mag_int_a_reg2);
	altbarrel_shift3 :  FloatConv_altbarrel_shift_lof
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_altbarrel_shift3_data,
		distance => leading_zeroes,
		result => wire_altbarrel_shift3_result
	  );
	altpriority_encoder2 :  FloatConv_altpriority_encoder_0c6
	  PORT MAP ( 
		data => prio_mag_int_a,
		q => wire_altpriority_encoder2_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_cout_reg <= wire_add_sub4_cout;
			END IF;
		END IF;
	END PROCESS;
	loop57 : FOR i IN 0 TO 26 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_w_lg_q69w70w(i) <= wire_add_1_adder1_cout_reg_w_lg_q69w(0) AND wire_mantissa_pre_round_reg_w_q_range68w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 26 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_q67w(i) <= add_1_adder1_cout_reg AND add_1_adder2_reg(i);
	END GENERATE loop58;
	wire_add_1_adder1_cout_reg_w_lg_q69w(0) <= NOT add_1_adder1_cout_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_reg <= wire_add_sub4_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_cout_reg <= wire_add_sub5_cout;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_reg <= wire_add_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_reg <= add_1_w;
			END IF;
		END IF;
	END PROCESS;
	loop59 : FOR i IN 0 TO 52 GENERATE 
		wire_add_1_reg_w_lg_w_lg_q76w77w(i) <= wire_add_1_reg_w_lg_q76w(0) AND mantissa_pre_round_reg(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 52 GENERATE 
		wire_add_1_reg_w_lg_q75w(i) <= add_1_reg AND mantissa_post_round(i);
	END GENERATE loop60;
	wire_add_1_reg_w_lg_q76w(0) <= NOT add_1_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg <= exponent_bus_pre_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg2 <= exponent_bus_pre_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg3 <= exponent_bus_pre;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg <= mag_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg2 <= mag_int_a_reg;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_pre_round_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_pre_round_reg <= mantissa_pre_round;
			END IF;
		END IF;
	END PROCESS;
	wire_mantissa_pre_round_reg_w_q_range68w <= mantissa_pre_round_reg(52 DOWNTO 26);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN priority_encoder_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN priority_encoder_reg <= wire_altpriority_encoder2_q;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_reg <= result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg1 <= sign_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg2 <= sign_int_a_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg3 <= sign_int_a_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg4 <= sign_int_a_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg5 <= sign_int_a_reg4;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_datab <= "000000000000000000000000000000000000000000000000000000000000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 63,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => invert_int_a,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	wire_add_sub4_datab <= "00000000000000000000000001";
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 26,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub4_cout,
		dataa => mantissa_pre_round(25 DOWNTO 0),
		datab => wire_add_sub4_datab,
		result => wire_add_sub4_result
	  );
	wire_add_sub5_datab <= "000000000000000000000000001";
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 27,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub5_cout,
		dataa => mantissa_pre_round(52 DOWNTO 26),
		datab => wire_add_sub5_datab,
		result => wire_add_sub5_result
	  );
	wire_add_sub6_datab <= "00000000001";
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 11,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_bus_pre_reg,
		datab => wire_add_sub6_datab,
		result => wire_add_sub6_result
	  );
	exponent_value :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 11,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => const_bias_value_add_width_int_w,
		datab => minus_leading_zero,
		result => wire_exponent_value_result
	  );
	loop61 : FOR i IN 0 TO 10 GENERATE 
		wire_below_bias_value_w_lg_w_lg_alb21w22w(i) <= wire_below_bias_value_w_lg_alb21w(0) AND exponent_output_w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 10 GENERATE 
		wire_below_bias_value_w_lg_alb20w(i) <= wire_below_bias_value_alb AND exceptions_value(i);
	END GENERATE loop62;
	wire_below_bias_value_w_lg_alb21w(0) <= NOT wire_below_bias_value_alb;
	below_bias_value :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		alb => wire_below_bias_value_alb,
		dataa => exponent_output_w,
		datab => bias_value_w
	  );

 END RTL; --FloatConv_altfp_convert_2gn
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FloatConv IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END FloatConv;


ARCHITECTURE RTL OF floatconv IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (63 DOWNTO 0);



	COMPONENT FloatConv_altfp_convert_2gn
	PORT (
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(63 DOWNTO 0);

	FloatConv_altfp_convert_2gn_component : FloatConv_altfp_convert_2gn
	PORT MAP (
		aclr => aclr,
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "FIXED2FLOAT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "64"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "11"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "12"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "52"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "64"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 64 0 INPUT NODEFVAL "dataa[63..0]"
-- Retrieval info: CONNECT: @dataa 0 0 64 0 dataa 0 0 64 0
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL FloatConv.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FloatConv.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FloatConv.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FloatConv_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FloatConv.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FloatConv.cmp TRUE TRUE
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX NUMERIC "1"
-- Retrieval info: LIB_FILE: lpm
