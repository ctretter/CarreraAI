-- AvalonSPI.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AvalonSPI is
	port (
		stsinkvalid   : in    std_logic                    := '0';             --   avalon_streaming_sink.valid
		stsinkdata    : in    std_logic_vector(7 downto 0) := (others => '0'); --                        .data
		stsinkready   : out   std_logic;                                       --                        .ready
		stsourceready : in    std_logic                    := '0';             -- avalon_streaming_source.ready
		stsourcevalid : out   std_logic;                                       --                        .valid
		stsourcedata  : out   std_logic_vector(7 downto 0);                    --                        .data
		sysclk        : in    std_logic                    := '0';             --              clock_sink.clk
		nreset        : in    std_logic                    := '0';             --        clock_sink_reset.reset_n
		mosi          : in    std_logic                    := '0';             --                export_0.mosi
		nss           : in    std_logic                    := '0';             --                        .nss
		miso          : inout std_logic                    := '0';             --                        .miso
		sclk          : in    std_logic                    := '0'              --                        .sclk
	);
end entity AvalonSPI;

architecture rtl of AvalonSPI is
	component SPIPhy is
		generic (
			SYNC_DEPTH : integer := 2
		);
		port (
			sysclk        : in    std_logic                    := 'X';             -- clk
			nreset        : in    std_logic                    := 'X';             -- reset_n
			mosi          : in    std_logic                    := 'X';             -- export
			nss           : in    std_logic                    := 'X';             -- export
			miso          : inout std_logic                    := 'X';             -- export
			sclk          : in    std_logic                    := 'X';             -- export
			stsourceready : in    std_logic                    := 'X';             -- ready
			stsourcevalid : out   std_logic;                                       -- valid
			stsourcedata  : out   std_logic_vector(7 downto 0);                    -- data
			stsinkvalid   : in    std_logic                    := 'X';             -- valid
			stsinkdata    : in    std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stsinkready   : out   std_logic                                        -- ready
		);
	end component SPIPhy;

begin

	spislave_0 : component SPIPhy
		generic map (
			SYNC_DEPTH => 2
		)
		port map (
			sysclk        => sysclk,        --              clock_sink.clk
			nreset        => nreset,        --        clock_sink_reset.reset_n
			mosi          => mosi,          --                export_0.export
			nss           => nss,           --                        .export
			miso          => miso,          --                        .export
			sclk          => sclk,          --                        .export
			stsourceready => stsourceready, -- avalon_streaming_source.ready
			stsourcevalid => stsourcevalid, --                        .valid
			stsourcedata  => stsourcedata,  --                        .data
			stsinkvalid   => stsinkvalid,   --   avalon_streaming_sink.valid
			stsinkdata    => stsinkdata,    --                        .data
			stsinkready   => stsinkready    --                        .ready
		);

end architecture rtl; -- of AvalonSPI
