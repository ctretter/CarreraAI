-------------------------------------------------------------------------------
-- Title      : Testbench for design "PwrOnReset"
-- Project    : 
-------------------------------------------------------------------------------
-- $Id: tbPwrOnReset-e.vhd 3 2011-09-10 08:35:02Z mroland $
-------------------------------------------------------------------------------
-- Author     : Copyright 2003: Markus Pfaff
-- Standard   : Using VHDL'93
-- Simulation : Model Technology Modelsim
-- Synthesis  : Exemplar Leonardo
-------------------------------------------------------------------------------
-- Description:
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

use work.Global.all;

-----------------------------------------------------------------------------------------

entity tbPwrOnReset is

end entity tbPwrOnReset;

