-------------------------------------------------------------------------------
-- Title      : Testbench for design "Oscillator"
-- Project    : IP
-------------------------------------------------------------------------------
-- $Id: tbOscillator-e.vhd 3 2011-09-10 08:35:02Z mroland $
-------------------------------------------------------------------------------
-- Author     : Copyright 2003: Markus Pfaff
-- Standard   : Using VHDL'93
-- Simulation : Model Technology Modelsim
-- Synthesis  : Exemplar Leonardo
-------------------------------------------------------------------------------
-- Description:
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity tbOscillator is

end entity tbOscillator;

