------------------------------------------------------------
--author: tretterch
--date:	  03-15-2017
--Descr.: Interface of cordic implementation for 
--	  exponential function
------------------------------------------------------------
--Rev	 author		date		comment
--0.1	tretterch     03-15-2017      initial implementation
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all
use ieee.numeric_std.all;
use ieee.fixed_generic_pkg.all;
use ieee.fixed_pkg.all

entity Cordic is
	generic();
	port(
		
	    );
end Cordic
