Exponential_inst : Exponential PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
